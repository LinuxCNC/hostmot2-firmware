library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from usb.obj
-- On 8/ 3/2009

entity usbrom is
	port (
	addr: in std_logic_vector(10 downto 0);
	clk: in std_logic;
	din: in std_logic_vector(15 downto 0);
	dout: out std_logic_vector(15 downto 0);
	we: in std_logic);
end usbrom;

architecture syn of usbrom is
   type ram_type is array (0 to 2047) of std_logic_vector(15 downto 0);
   signal RAM : ram_type := 
   (
   x"0000", x"0000", x"6433", x"0100", x"E7E3", x"203E", x"0000", x"0000",
   x"0000", x"0101", x"B07B", x"0100", x"B7E3", x"0100", x"B7E6", x"0109",
   x"B7E7", x"013D", x"B7E8", x"0100", x"B7E9", x"0101", x"B07B", x"707B",
   x"97CD", x"A7C7", x"3031", x"0100", x"B07B", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"707C", x"B7D2", x"0101", x"B07B", x"77D2", x"C416",
   x"B416", x"0100", x"B7E6", x"0109", x"B7E7", x"013D", x"B7E8", x"0100",
   x"B7E9", x"77E6", x"E7C7", x"B7E6", x"77E7", x"F7C6", x"B7E7", x"77E8",
   x"F7C6", x"B7E8", x"77E9", x"F7C6", x"B7E9", x"4015", x"6433", x"0100",
   x"B07A", x"01EE", x"E06F", x"2047", x"0000", x"01FF", x"B7F7", x"0150",
   x"0800", x"0104", x"0A00", x"0100", x"B7F3", x"0100", x"B416", x"0100",
   x"B417", x"0100", x"B7D5", x"63CD", x"77D2", x"B7CF", x"01C0", x"A7D2",
   x"304D", x"0000", x"01FF", x"B7F3", x"011F", x"A7CF", x"B7E0", x"01C0",
   x"A7CF", x"B7DF", x"0000", x"0000", x"01C0", x"E7DF", x"206F", x"0000",
   x"0000", x"01FF", x"E7CF", x"206F", x"0000", x"0000", x"1047", x"0180",
   x"E7DF", x"208E", x"013F", x"A7CF", x"B7E1", x"01FF", x"B7D5", x"0000",
   x"77E1", x"C7C6", x"0200", x"0200", x"0200", x"0200", x"0200", x"0B00",
   x"0300", x"A7D6", x"0900", x"0700", x"A7D7", x"C7D8", x"0B00", x"0000",
   x"0000", x"7900", x"B7CF", x"0D01", x"0000", x"0000", x"77CF", x"B800",
   x"0C01", x"01C0", x"A7CF", x"B7DF", x"01F0", x"A7CF", x"B7F6", x"013F",
   x"A7CF", x"B7E1", x"0108", x"A7CF", x"B7EA", x"0104", x"A7CF", x"B7D0",
   x"0103", x"A7CF", x"B7D1", x"0120", x"A7CF", x"B7CE", x"0150", x"E7F6",
   x"3127", x"0000", x"0000", x"01C0", x"E7DF", x"20BB", x"0120", x"E7CE",
   x"20BB", x"0100", x"E7D5", x"30BA", x"0000", x"0000", x"7900", x"B800",
   x"0C01", x"10BB", x"6397", x"0140", x"E7DF", x"2127", x"0104", x"E7D0",
   x"20CF", x"0100", x"E7D5", x"30CD", x"0000", x"0000", x"7900", x"B800",
   x"7901", x"B801", x"0C02", x"0D02", x"10CF", x"6397", x"6397", x"0120",
   x"E7CE", x"2127", x"0100", x"E7D1", x"20DF", x"0110", x"A7CF", x"30DE",
   x"0000", x"7900", x"B800", x"0C01", x"0D01", x"10DF", x"6397", x"0101",
   x"E7D1", x"20EF", x"0110", x"A7CF", x"30ED", x"0000", x"7900", x"B800",
   x"7901", x"B801", x"0C02", x"0D02", x"10EF", x"6397", x"6397", x"0102",
   x"E7D1", x"2105", x"0110", x"A7CF", x"3101", x"0000", x"7900", x"B800",
   x"7901", x"B801", x"7902", x"B802", x"7903", x"B803", x"0C04", x"0D04",
   x"1105", x"6397", x"6397", x"6397", x"6397", x"0103", x"E7D1", x"2127",
   x"0110", x"A7CF", x"311F", x"0000", x"7900", x"B800", x"7901", x"B801",
   x"7902", x"B802", x"7903", x"B803", x"7904", x"B804", x"7905", x"B805",
   x"7906", x"B806", x"7907", x"B807", x"0C08", x"0D08", x"1127", x"6397",
   x"6397", x"6397", x"6397", x"6397", x"6397", x"6397", x"6397", x"0100",
   x"E7D5", x"212D", x"0000", x"0100", x"B7CF", x"0100", x"B800", x"0100",
   x"E7D5", x"3143", x"0000", x"7900", x"B7CF", x"0D01", x"B800", x"0C01",
   x"0400", x"E7D3", x"0600", x"F7D4", x"5143", x"0000", x"0000", x"0110",
   x"8411", x"B411", x"1047", x"77CF", x"2091", x"0000", x"0100", x"B7D5",
   x"0100", x"B800", x"0150", x"0800", x"0104", x"0A00", x"0000", x"0000",
   x"7800", x"B7CF", x"0C01", x"0000", x"0000", x"01C0", x"A7CF", x"B7DF",
   x"01F0", x"A7CF", x"B7F6", x"0108", x"A7CF", x"B7EA", x"0104", x"A7CF",
   x"B7D0", x"0103", x"A7CF", x"B7D1", x"0120", x"A7CF", x"B7CE", x"01C0",
   x"E7DF", x"2258", x"011F", x"A7CF", x"B7E0", x"0120", x"A7CF", x"B7CE",
   x"0500", x"B7DB", x"0700", x"B7DC", x"010F", x"E7E0", x"5190", x"0000",
   x"0000", x"0110", x"0900", x"0104", x"0B00", x"0500", x"C7E0", x"0900",
   x"0700", x"D7C6", x"0B00", x"0120", x"E7CE", x"218C", x"0000", x"0000",
   x"7800", x"0C01", x"B900", x"118F", x"0000", x"7900", x"6401", x"1254",
   x"0120", x"E7CE", x"21F2", x"0000", x"0000", x"01F7", x"E7CF", x"219D",
   x"0000", x"7800", x"0C01", x"B07A", x"11F1", x"01F8", x"E7CF", x"21AF",
   x"0100", x"E41A", x"21AA", x"0000", x"0000", x"0000", x"7800", x"0C01",
   x"B7D9", x"11AE", x"0000", x"7800", x"0C01", x"B7DD", x"11F1", x"01F9",
   x"E7CF", x"21C1", x"0100", x"E41A", x"21BC", x"0000", x"0000", x"0000",
   x"7800", x"0C01", x"B7DA", x"11C0", x"0000", x"7800", x"0C01", x"B7DE",
   x"11F1", x"01FA", x"E7CF", x"21D9", x"0100", x"E41A", x"21D0", x"0000",
   x"7800", x"0C01", x"C7D9", x"B7D9", x"77DA", x"D7C6", x"B7DA", x"11D8",
   x"0000", x"7800", x"0C01", x"C7DD", x"B7DD", x"77DE", x"D7C6", x"B7DE",
   x"11F1", x"01FD", x"E7CF", x"21E1", x"0000", x"7800", x"0C01", x"B7F0",
   x"11F1", x"01FE", x"E7CF", x"21F1", x"0000", x"7800", x"0C01", x"B7D2",
   x"0000", x"0000", x"015A", x"E7D2", x"21F0", x"0000", x"0000", x"103E",
   x"11F1", x"1254", x"01D0", x"E7CF", x"21F9", x"0000", x"0137", x"6401",
   x"1254", x"01D1", x"E7CF", x"2200", x"0000", x"0149", x"6401", x"1254",
   x"01D2", x"E7CF", x"2207", x"0000", x"0134", x"6401", x"1254", x"01D3",
   x"E7CF", x"220E", x"0000", x"0133", x"6401", x"1254", x"01DA", x"E7CF",
   x"2215", x"0000", x"0106", x"6401", x"1254", x"01DB", x"E7CF", x"221C",
   x"0000", x"742B", x"6401", x"1254", x"01DD", x"E7CF", x"2223", x"0000",
   x"0100", x"6401", x"1254", x"01DE", x"E7CF", x"222A", x"0000", x"0104",
   x"6401", x"1254", x"01DC", x"E7CF", x"2231", x"0000", x"0110", x"6401",
   x"1254", x"01D8", x"E7CF", x"223F", x"0000", x"0100", x"E41A", x"223C",
   x"0000", x"0000", x"77D9", x"123D", x"77DD", x"6401", x"1254", x"01D9",
   x"E7CF", x"224D", x"0000", x"0100", x"E41A", x"224A", x"0000", x"0000",
   x"77DA", x"124B", x"77DE", x"6401", x"1254", x"01DF", x"E7CF", x"2254",
   x"0000", x"015A", x"6401", x"1254", x"77DB", x"0900", x"77DC", x"0B00",
   x"013F", x"A7CF", x"B7E1", x"0150", x"E7F6", x"22BF", x"0107", x"A7CF",
   x"B7F6", x"0100", x"B7F4", x"0100", x"B7F5", x"0100", x"E7F6", x"226D",
   x"0101", x"B7F4", x"0100", x"B7F5", x"129D", x"0101", x"E7F6", x"2275",
   x"0102", x"B7F4", x"01FF", x"B7F5", x"129D", x"0102", x"E7F6", x"227D",
   x"0104", x"B7F4", x"0100", x"B7F5", x"129D", x"0103", x"E7F6", x"2285",
   x"0108", x"B7F4", x"01FF", x"B7F5", x"129D", x"0104", x"E7F6", x"228D",
   x"0110", x"B7F4", x"01FF", x"B7F5", x"129D", x"0106", x"E7F6", x"2295",
   x"0140", x"B7F4", x"01FF", x"B7F5", x"129D", x"0107", x"E7F6", x"229D",
   x"0180", x"B7F4", x"01FF", x"B7F5", x"129D", x"01D0", x"B7F0", x"0118",
   x"B7F1", x"741B", x"B7F2", x"77F0", x"E7C7", x"B7F0", x"77F1", x"F7C6",
   x"B7F1", x"42B8", x"0000", x"0000", x"01D0", x"B7F0", x"0118", x"B7F1",
   x"77F2", x"E7C7", x"B7F2", x"42B8", x"0180", x"8411", x"B411", x"1047",
   x"7089", x"97F5", x"A7F4", x"32A3", x"0000", x"0000", x"1390", x"0140",
   x"E7DF", x"2390", x"0104", x"E7D0", x"22D5", x"0100", x"E41A", x"22CF",
   x"0000", x"7800", x"B7D9", x"7801", x"B7DA", x"0C02", x"12D5", x"0000",
   x"7800", x"B7DD", x"7801", x"B7DE", x"0C02", x"0100", x"E41A", x"22EE",
   x"0000", x"0000", x"77F7", x"22E2", x"0000", x"77D9", x"0900", x"77DA",
   x"0B00", x"12ED", x"77D9", x"B068", x"A7C9", x"B7CB", x"77DA", x"B069",
   x"0100", x"0B00", x"0160", x"C7CB", x"0900", x"12F3", x"77DD", x"0900",
   x"77DE", x"C7D8", x"0B00", x"0100", x"E41A", x"22FF", x"0000", x"0000",
   x"77F7", x"22FE", x"01FF", x"E7D9", x"0103", x"F7DA", x"1303", x"01FF",
   x"E7DD", x"0103", x"F7DE", x"430D", x"0000", x"0000", x"0100", x"0900",
   x"0104", x"0B00", x"0120", x"8411", x"B411", x"0120", x"E7CE", x"2350",
   x"0100", x"E7D1", x"2319", x"0000", x"7800", x"B900", x"0C01", x"77C7",
   x"6411", x"0101", x"E7D1", x"2324", x"0000", x"7800", x"B900", x"7801",
   x"B901", x"0C02", x"77C8", x"6411", x"0102", x"E7D1", x"2333", x"0000",
   x"7800", x"B900", x"7801", x"B901", x"7802", x"B902", x"7803", x"B903",
   x"0C04", x"77CA", x"6411", x"0103", x"E7D1", x"234A", x"0000", x"7800",
   x"B900", x"7801", x"B901", x"7802", x"B902", x"7803", x"B903", x"7804",
   x"B904", x"7805", x"B905", x"7806", x"B906", x"7807", x"B907", x"0C08",
   x"77CC", x"6411", x"77F7", x"334F", x"0000", x"0000", x"B06E", x"1390",
   x"77F7", x"3355", x"0000", x"0000", x"B06D", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0100", x"E7D1", x"2362", x"0000", x"7900", x"6401",
   x"77C7", x"6411", x"0101", x"E7D1", x"236C", x"0000", x"7900", x"6401",
   x"7901", x"6401", x"77C8", x"6411", x"0102", x"E7D1", x"237A", x"0000",
   x"7900", x"6401", x"7901", x"6401", x"7902", x"6401", x"7903", x"6401",
   x"77CA", x"6411", x"0103", x"E7D1", x"2390", x"0000", x"7900", x"6401",
   x"7901", x"6401", x"7902", x"6401", x"7903", x"6401", x"7904", x"6401",
   x"7905", x"6401", x"7906", x"6401", x"7907", x"6401", x"77CC", x"6411",
   x"7800", x"2150", x"0000", x"0000", x"1047", x"0000", x"0000", x"01D0",
   x"B7F0", x"0118", x"B7F1", x"741B", x"B7F2", x"77F0", x"E7C7", x"B7F0",
   x"77F1", x"F7C6", x"B7F1", x"43B4", x"0000", x"01D0", x"B7F0", x"0118",
   x"B7F1", x"77F2", x"E7C7", x"B7F2", x"43B4", x"0000", x"77F3", x"33B4",
   x"0140", x"8411", x"B411", x"1047", x"0101", x"B07B", x"707B", x"97CD",
   x"A7C7", x"339D", x"0000", x"0100", x"B07B", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"707C", x"B7D2", x"0101", x"B07B", x"77D2", x"C416",
   x"B416", x"77D2", x"B800", x"0C01", x"1800", x"01D0", x"B7F0", x"0118",
   x"B7F1", x"741B", x"B7F2", x"77F0", x"E7C7", x"B7F0", x"77F1", x"F7C6",
   x"B7F1", x"43EA", x"0000", x"01D0", x"B7F0", x"0118", x"B7F1", x"77F2",
   x"E7C7", x"B7F2", x"43EA", x"0000", x"77F3", x"33EA", x"0140", x"8411",
   x"B411", x"1047", x"0101", x"B07B", x"707B", x"97CD", x"A7C7", x"33D3",
   x"0000", x"0100", x"B07B", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"707C", x"B7D2", x"0101", x"B07B", x"77D2", x"C416", x"B416", x"0000",
   x"1800", x"B7D2", x"707B", x"97CD", x"A7C8", x"3402", x"0105", x"B07B",
   x"0107", x"B07B", x"77D2", x"B07C", x"C417", x"B417", x"0101", x"B07B",
   x"1800", x"B7EB", x"77EA", x"3800", x"0500", x"C7EB", x"0900", x"0700",
   x"D7C6", x"0B00", x"0100", x"E41A", x"242D", x"0000", x"0000", x"77F7",
   x"3428", x"77D9", x"C7EB", x"B7D9", x"77DA", x"D7C6", x"B7DA", x"142C",
   x"0500", x"B7D9", x"0700", x"B7DA", x"1432", x"0500", x"B7DD", x"0700",
   x"E7D8", x"B7DE", x"1800", x"0100", x"B7D2", x"B410", x"B411", x"B412",
   x"B413", x"B415", x"B416", x"B417", x"B418", x"B419", x"B41A", x"B42B",
   x"B7F0", x"B7C6", x"0101", x"B7C7", x"0102", x"B7C8", x"0103", x"B7C9",
   x"0104", x"B7CA", x"0108", x"B7CC", x"01FF", x"B7CD", x"B41B", x"01F0",
   x"B7D6", x"0103", x"B7D7", x"010C", x"B7D8", x"01C0", x"B7DF", x"017A",
   x"B7D9", x"0100", x"B7DA", x"0100", x"B7DD", x"0100", x"B7DE", x"01B4",
   x"B7D3", x"0107", x"B7D4", x"1800", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000"
);

signal daddr: std_logic_vector(10 downto 0);

begin
   ausbrom: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (we = '1') then
            RAM(conv_integer(addr)) <= din;
         end if;
         daddr <= addr;
      end if; -- clk 
   end process;

   dout <= RAM(conv_integer(daddr));
end;
