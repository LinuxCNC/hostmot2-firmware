library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from testrom.bin
-- On 1/ 5/2009

entity testrom is
	port (
	addr: in std_logic_vector(10 downto 0);
	clk: in std_logic;
	din: in std_logic_vector(23 downto 0);
	dout: out std_logic_vector(23 downto 0);
	we: in std_logic);
end testrom;

architecture syn of testrom is
   type ram_type is array (0 to 2047) of std_logic_vector(23 downto 0);
   signal RAM : ram_type := 
   (
   x"000000", x"000000", x"012710", x"B00003", x"010000",
   x"B00004", x"02FFFF", x"03FFFF", x"B00007", x"010005",
   x"B00004", x"020000", x"03FFFB", x"A00004", x"B00000",
   x"200009", x"400001", x"600007", x"030000", x"32001B",
   x"400005", x"C00003", x"B00005", x"400000", x"D00004",
   x"B00000", x"200021", x"400005", x"E00003", x"B00005",
   x"400000", x"F00004", x"B00000", x"200010", x"000000",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF",
   x"FFFFFF", x"FFFFFF", x"01ABCD");

signal daddr: std_logic_vector(10 downto 0);

begin
   atestrom: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (we = '1') then
            RAM(conv_integer(addr)) <= din;
         end if;
         daddr <= addr;
      end if; -- clk 
   end process;

   dout <= RAM(conv_integer(daddr));
end;
