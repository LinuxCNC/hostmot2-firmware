library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from usb.obj
-- On11/ 9/2009

entity usbrom is
	port (
	addr: in std_logic_vector(9 downto 0);
	clk: in std_logic;
	din: in std_logic_vector(15 downto 0);
	dout: out std_logic_vector(15 downto 0);
	we: in std_logic);
end usbrom;

architecture syn of usbrom is
   type ram_type is array (0 to 1023) of std_logic_vector(15 downto 0);
   signal RAM : ram_type := 
   (
   x"0000", x"0000", x"63C7", x"0100", x"E7E3", x"203C", x"0000", x"0000",
   x"0000", x"0101", x"B07B", x"0100", x"B7E3", x"0100", x"B7E6", x"0109",
   x"B7E7", x"013D", x"B7E8", x"0100", x"B7E9", x"0101", x"B07B", x"707B",
   x"97CD", x"A7C7", x"302F", x"0100", x"B07B", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"707C", x"B7D2", x"0101", x"B07B", x"77D2", x"0100",
   x"B7E6", x"0109", x"B7E7", x"013D", x"B7E8", x"0100", x"B7E9", x"77E6",
   x"E7C7", x"B7E6", x"77E7", x"F7C6", x"B7E7", x"77E8", x"F7C6", x"B7E8",
   x"77E9", x"F7C6", x"B7E9", x"4015", x"63C7", x"0100", x"B07A", x"01EE",
   x"E06F", x"2045", x"0000", x"01FF", x"B7F7", x"0150", x"0800", x"0104",
   x"0A00", x"0100", x"B7F3", x"0100", x"B7F6", x"0100", x"B7D5", x"6363",
   x"77D2", x"B7CF", x"01C0", x"A7D2", x"304B", x"0000", x"01FF", x"B7F3",
   x"011F", x"A7CF", x"B7E0", x"01C0", x"A7CF", x"B7DF", x"0000", x"0000",
   x"01C0", x"E7DF", x"206B", x"0000", x"0000", x"01FF", x"E7CF", x"206B",
   x"0000", x"0000", x"1045", x"0180", x"E7DF", x"208A", x"013F", x"A7CF",
   x"B7E1", x"01FF", x"B7D5", x"0000", x"77E1", x"C7C6", x"0200", x"0200",
   x"0200", x"0200", x"0200", x"0B00", x"0300", x"A7D6", x"0900", x"0700",
   x"A7D7", x"C7D8", x"0B00", x"0000", x"0000", x"7900", x"B7CF", x"0D01",
   x"0000", x"0000", x"77CF", x"B800", x"0C01", x"01C0", x"A7CF", x"B7DF",
   x"013F", x"A7CF", x"B7E1", x"0108", x"A7CF", x"B7EA", x"0104", x"A7CF",
   x"B7D0", x"0103", x"A7CF", x"B7D1", x"0120", x"A7CF", x"B7CE", x"01C0",
   x"E7DF", x"20AF", x"0120", x"E7CE", x"20AF", x"0100", x"E7D5", x"30AE",
   x"0000", x"0000", x"7900", x"B800", x"0C01", x"10AF", x"632F", x"0140",
   x"E7DF", x"211B", x"0104", x"E7D0", x"20C3", x"0100", x"E7D5", x"30C1",
   x"0000", x"0000", x"7900", x"B800", x"7901", x"B801", x"0C02", x"0D02",
   x"10C3", x"632F", x"632F", x"0120", x"E7CE", x"211B", x"0100", x"E7D1",
   x"20D3", x"0110", x"A7CF", x"30D2", x"0000", x"7900", x"B800", x"0C01",
   x"0D01", x"10D3", x"632F", x"0101", x"E7D1", x"20E3", x"0110", x"A7CF",
   x"30E1", x"0000", x"7900", x"B800", x"7901", x"B801", x"0C02", x"0D02",
   x"10E3", x"632F", x"632F", x"0102", x"E7D1", x"20F9", x"0110", x"A7CF",
   x"30F5", x"0000", x"7900", x"B800", x"7901", x"B801", x"7902", x"B802",
   x"7903", x"B803", x"0C04", x"0D04", x"10F9", x"632F", x"632F", x"632F",
   x"632F", x"0103", x"E7D1", x"211B", x"0110", x"A7CF", x"3113", x"0000",
   x"7900", x"B800", x"7901", x"B801", x"7902", x"B802", x"7903", x"B803",
   x"7904", x"B804", x"7905", x"B805", x"7906", x"B806", x"7907", x"B807",
   x"0C08", x"0D08", x"111B", x"632F", x"632F", x"632F", x"632F", x"632F",
   x"632F", x"632F", x"632F", x"0100", x"E7D5", x"2121", x"0000", x"0100",
   x"B7CF", x"0100", x"B800", x"0100", x"E7D5", x"3137", x"0000", x"7900",
   x"B7CF", x"0D01", x"B800", x"0C01", x"0400", x"E7D3", x"0600", x"F7D4",
   x"5137", x"0000", x"0000", x"0110", x"8411", x"B411", x"1045", x"77CF",
   x"208D", x"0000", x"0100", x"B7D5", x"0100", x"B800", x"0100", x"B7F3",
   x"0150", x"0800", x"0104", x"0A00", x"0000", x"0000", x"0100", x"B7F6",
   x"7800", x"B7CF", x"0C01", x"0000", x"0000", x"01C0", x"A7CF", x"B7DF",
   x"0108", x"A7CF", x"B7EA", x"0104", x"A7CF", x"B7D0", x"0103", x"A7CF",
   x"B7D1", x"0120", x"A7CF", x"B7CE", x"01C0", x"E7DF", x"2254", x"011F",
   x"A7CF", x"B7E0", x"0120", x"A7CF", x"B7CE", x"0500", x"B7DB", x"0700",
   x"B7DC", x"010F", x"E7E0", x"5185", x"0000", x"0000", x"0110", x"0900",
   x"0104", x"0B00", x"0500", x"C7E0", x"0900", x"0700", x"D7C6", x"0B00",
   x"0120", x"E7CE", x"2181", x"0000", x"0000", x"7800", x"0C01", x"B900",
   x"1184", x"0000", x"7900", x"6395", x"1250", x"0120", x"E7CE", x"21E7",
   x"0000", x"0000", x"01F7", x"E7CF", x"2192", x"0000", x"7800", x"0C01",
   x"B07A", x"11E6", x"01F8", x"E7CF", x"21A4", x"0100", x"E41A", x"219F",
   x"0000", x"0000", x"0000", x"7800", x"0C01", x"B7D9", x"11A3", x"0000",
   x"7800", x"0C01", x"B7DD", x"11E6", x"01F9", x"E7CF", x"21B6", x"0100",
   x"E41A", x"21B1", x"0000", x"0000", x"0000", x"7800", x"0C01", x"B7DA",
   x"11B5", x"0000", x"7800", x"0C01", x"B7DE", x"11E6", x"01FA", x"E7CF",
   x"21CE", x"0100", x"E41A", x"21C5", x"0000", x"7800", x"0C01", x"C7D9",
   x"B7D9", x"77DA", x"D7C6", x"B7DA", x"11CD", x"0000", x"7800", x"0C01",
   x"C7DD", x"B7DD", x"77DE", x"D7C6", x"B7DE", x"11E6", x"01FD", x"E7CF",
   x"21D6", x"0000", x"7800", x"0C01", x"B7F0", x"11E6", x"01FE", x"E7CF",
   x"21E6", x"0000", x"7800", x"0C01", x"B7D2", x"0000", x"0000", x"015A",
   x"E7D2", x"21E5", x"0000", x"0000", x"103C", x"11E6", x"1250", x"01D0",
   x"E7CF", x"21EE", x"0000", x"0137", x"6395", x"1250", x"01D1", x"E7CF",
   x"21F5", x"0000", x"0149", x"6395", x"1250", x"01D2", x"E7CF", x"21FC",
   x"0000", x"0134", x"6395", x"1250", x"01D3", x"E7CF", x"2203", x"0000",
   x"0133", x"6395", x"1250", x"01D4", x"E7CF", x"220A", x"0000", x"0100",
   x"6395", x"1250", x"01DA", x"E7CF", x"2211", x"0000", x"0105", x"6395",
   x"1250", x"01DB", x"E7CF", x"2218", x"0000", x"742B", x"6395", x"1250",
   x"01DD", x"E7CF", x"221F", x"0000", x"0100", x"6395", x"1250", x"01DE",
   x"E7CF", x"2226", x"0000", x"0104", x"6395", x"1250", x"01DC", x"E7CF",
   x"222D", x"0000", x"0110", x"6395", x"1250", x"01D8", x"E7CF", x"223B",
   x"0000", x"0100", x"E41A", x"2238", x"0000", x"0000", x"77D9", x"1239",
   x"77DD", x"6395", x"1250", x"01D9", x"E7CF", x"2249", x"0000", x"0100",
   x"E41A", x"2246", x"0000", x"0000", x"77DA", x"1247", x"77DE", x"6395",
   x"1250", x"01DF", x"E7CF", x"2250", x"0000", x"015A", x"6395", x"1250",
   x"77DB", x"0900", x"77DC", x"0B00", x"013F", x"A7CF", x"B7E1", x"0140",
   x"E7DF", x"2328", x"0104", x"E7D0", x"226D", x"0100", x"E41A", x"2267",
   x"0000", x"7800", x"B7D9", x"7801", x"B7DA", x"0C02", x"126D", x"0000",
   x"7800", x"B7DD", x"7801", x"B7DE", x"0C02", x"0100", x"E41A", x"2286",
   x"0000", x"0000", x"77F7", x"227A", x"0000", x"77D9", x"0900", x"77DA",
   x"0B00", x"1285", x"77D9", x"B068", x"A7C9", x"B7CB", x"77DA", x"B069",
   x"0100", x"0B00", x"0160", x"C7CB", x"0900", x"128B", x"77DD", x"0900",
   x"77DE", x"C7D8", x"0B00", x"0100", x"E41A", x"2297", x"0000", x"0000",
   x"77F7", x"2296", x"01FF", x"E7D9", x"0103", x"F7DA", x"129B", x"01FF",
   x"E7DD", x"0103", x"F7DE", x"42A5", x"0000", x"0000", x"0100", x"0900",
   x"0104", x"0B00", x"0120", x"8411", x"B411", x"0120", x"E7CE", x"22E8",
   x"0100", x"E7D1", x"22B1", x"0000", x"7800", x"B900", x"0C01", x"77C7",
   x"63A5", x"0101", x"E7D1", x"22BC", x"0000", x"7800", x"B900", x"7801",
   x"B901", x"0C02", x"77C8", x"63A5", x"0102", x"E7D1", x"22CB", x"0000",
   x"7800", x"B900", x"7801", x"B901", x"7802", x"B902", x"7803", x"B903",
   x"0C04", x"77CA", x"63A5", x"0103", x"E7D1", x"22E2", x"0000", x"7800",
   x"B900", x"7801", x"B901", x"7802", x"B902", x"7803", x"B903", x"7804",
   x"B904", x"7805", x"B905", x"7806", x"B906", x"7807", x"B907", x"0C08",
   x"77CC", x"63A5", x"77F7", x"32E7", x"0000", x"0000", x"B06E", x"1328",
   x"77F7", x"32ED", x"0000", x"0000", x"B06D", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0100", x"E7D1", x"22FA", x"0000", x"7900", x"6395",
   x"77C7", x"63A5", x"0101", x"E7D1", x"2304", x"0000", x"7900", x"6395",
   x"7901", x"6395", x"77C8", x"63A5", x"0102", x"E7D1", x"2312", x"0000",
   x"7900", x"6395", x"7901", x"6395", x"7902", x"6395", x"7903", x"6395",
   x"77CA", x"63A5", x"0103", x"E7D1", x"2328", x"0000", x"7900", x"6395",
   x"7901", x"6395", x"7902", x"6395", x"7903", x"6395", x"7904", x"6395",
   x"7905", x"6395", x"7906", x"6395", x"7907", x"6395", x"77CC", x"63A5",
   x"7800", x"2146", x"0000", x"0000", x"1045", x"0000", x"0000", x"01D0",
   x"B7F0", x"0118", x"B7F1", x"741B", x"B7F2", x"77F0", x"E7C7", x"B7F0",
   x"77F1", x"F7C6", x"B7F1", x"434C", x"0000", x"01D0", x"B7F0", x"0118",
   x"B7F1", x"77F2", x"E7C7", x"B7F2", x"434C", x"0000", x"77F3", x"334C",
   x"0140", x"8411", x"B411", x"1045", x"0101", x"B07B", x"707B", x"97CD",
   x"A7C7", x"3335", x"0000", x"0100", x"B07B", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"707C", x"B7D2", x"0101", x"B07B", x"77D2", x"77D2",
   x"B800", x"0C01", x"1800", x"01D0", x"B7F0", x"0118", x"B7F1", x"741B",
   x"B7F2", x"77F0", x"E7C7", x"B7F0", x"77F1", x"F7C6", x"B7F1", x"4380",
   x"0000", x"01D0", x"B7F0", x"0118", x"B7F1", x"77F2", x"E7C7", x"B7F2",
   x"4380", x"0000", x"77F3", x"3380", x"0140", x"8411", x"B411", x"1045",
   x"0101", x"B07B", x"707B", x"97CD", x"A7C7", x"3369", x"0000", x"0100",
   x"B07B", x"0000", x"0000", x"0000", x"0000", x"0000", x"707C", x"B7D2",
   x"0101", x"B07B", x"77D2", x"0000", x"1800", x"B7D2", x"707B", x"97CD",
   x"A7C8", x"3396", x"0105", x"B07B", x"0107", x"B07B", x"77D2", x"B07C",
   x"0000", x"0000", x"0101", x"B07B", x"1800", x"B7EB", x"77EA", x"3800",
   x"0500", x"C7EB", x"0900", x"0700", x"D7C6", x"0B00", x"0100", x"E41A",
   x"23C1", x"0000", x"0000", x"77F7", x"33BC", x"77D9", x"C7EB", x"B7D9",
   x"77DA", x"D7C6", x"B7DA", x"13C0", x"0500", x"B7D9", x"0700", x"B7DA",
   x"13C6", x"0500", x"B7DD", x"0700", x"E7D8", x"B7DE", x"1800", x"0100",
   x"B7D2", x"B410", x"B411", x"B41A", x"B42B", x"B7F0", x"B7C6", x"0101",
   x"B7C7", x"0102", x"B7C8", x"0103", x"B7C9", x"0104", x"B7CA", x"0108",
   x"B7CC", x"01FF", x"B7CD", x"B41B", x"01F0", x"B7D6", x"0103", x"B7D7",
   x"010C", x"B7D8", x"01C0", x"B7DF", x"017A", x"B7D9", x"0100", x"B7DA",
   x"0100", x"B7DD", x"0100", x"B7DE", x"01B4", x"B7D3", x"0107", x"B7D4",
   x"1800", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000"
);

signal daddr: std_logic_vector(9 downto 0);

begin
   ausbrom: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (we = '1') then
            RAM(conv_integer(addr)) <= din;
         end if;
         daddr <= addr;
      end if; -- clk 
   end process;

   dout <= RAM(conv_integer(daddr));
end;
