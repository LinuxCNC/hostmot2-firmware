library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from etherhm2.bin
-- On 6/18/2014

entity etherhm2 is
	port (
	addr: in std_logic_vector(11 downto 0);
	clk: in std_logic;
	din: in std_logic_vector(23 downto 0);
	dout: out std_logic_vector(23 downto 0);
	we: in std_logic);
end etherhm2;

architecture syn of etherhm2 is
   type ram_type is array (0 to 4095) of std_logic_vector(23 downto 0);
   signal RAM : ram_type := 
   (
   x"000000", x"000000", x"000000", x"010000", x"8F0000",
   x"01FFFF", x"B0007B", x"B0007A", x"010064", x"100410",
   x"010000", x"B0007A", x"100237", x"100361", x"1003BF",
   x"1002F5", x"40013A", x"330000", x"40012C", x"330017",
   x"010000", x"B00079", x"200019", x"010001", x"B00079",
   x"4B0000", x"B0007A", x"4000AC", x"33001F", x"400031",
   x"330012", x"40007C", x"B00150", x"01017F", x"850000",
   x"10009E", x"320012", x"010180", x"850000", x"000000",
   x"000000", x"010800", x"060000", x"E90006", x"320046",
   x"010806", x"060000", x"E90006", x"320034", x"000000",
   x"000000", x"200012", x"4000A8", x"E90013", x"330012",
   x"4000A9", x"E90014", x"330012", x"0104B6", x"840000",
   x"010806", x"060000", x"B000B6", x"010040", x"B000B4",
   x"1003D9", x"10018A", x"100199", x"10010D", x"200012",
   x"4000A8", x"E9000F", x"330012", x"4000A9", x"E90010",
   x"330012", x"49000B", x"E0008F", x"70008D", x"320057",
   x"49000B", x"E00090", x"70008D", x"32006C", x"000000",
   x"000000", x"200012", x"010180", x"840000", x"4000AD",
   x"B000B4", x"010800", x"060000", x"B000B6", x"10018A",
   x"1001D5", x"1001F0", x"01FFF2", x"C080AD", x"014001",
   x"060000", x"B8000B", x"000000", x"4000AD", x"060000",
   x"B80008", x"10010D", x"200012", x"490012", x"E000D8",
   x"330012", x"490013", x"060000", x"E00088", x"0B0000",
   x"B000DC", x"0104CB", x"840000", x"010195", x"850000",
   x"40007C", x"B00151", x"200469", x"B000B4", x"320010",
   x"010001", x"C08134", x"0104B6", x"840000", x"010180",
   x"850000", x"010008", x"C080B4", x"010800", x"060000",
   x"B000B6", x"10018A", x"1001D5", x"1001F7", x"4000B4",
   x"060000", x"B80013", x"010014", x"C080B4", x"014011",
   x"060000", x"B8000B", x"4000B4", x"060000", x"B80008",
   x"01000E", x"C080B4", x"40007C", x"B00152", x"10010D",
   x"40007C", x"B00153", x"200010", x"B0003C", x"4000AC",
   x"3300B6", x"000000", x"01C092", x"100154", x"40009F",
   x"B0009E", x"01C092", x"100141", x"012000", x"70009F",
   x"3200F8", x"010000", x"B0009E", x"013090", x"100141",
   x"01309C", x"100154", x"01FF00", x"70009F", x"060000",
   x"B000AC", x"320102", x"000000", x"01FFFF", x"C080AC",
   x"01307C", x"100154", x"018000", x"70009F", x"3200FE",
   x"010017", x"70009F", x"3300FE", x"013C00", x"70009F",
   x"3300FE", x"000000", x"01C07E", x"100154", x"010FFF",
   x"70009F", x"B000AD", x"B000AE", x"3200FE", x"014000",
   x"B0009E", x"01C086", x"100141", x"010238", x"B0009E",
   x"01C082", x"100141", x"10016A", x"10016A", x"10016A",
   x"C00083", x"70008E", x"B000AE", x"E000B9", x"3C00FE",
   x"B00041", x"400045", x"000000", x"000000", x"000000",
   x"000000", x"400041", x"B90000", x"400045", x"000000",
   x"000000", x"000000", x"000000", x"400041", x"B90001",
   x"01FFFC", x"C080AE", x"890002", x"3300DD", x"000000",
   x"010230", x"B0009E", x"01C082", x"100141", x"012800",
   x"B0009E", x"013090", x"100141", x"010001", x"C08130",
   x"01FFFA", x"C080AD", x"B0003D", x"280000", x"010231",
   x"B0009E", x"01C082", x"100141", x"012800", x"B0009E",
   x"013090", x"100141", x"010008", x"50812C", x"010001",
   x"C08132", x"010000", x"B0003D", x"280000", x"B0003E",
   x"4000B4", x"C00083", x"70008E", x"B000B5", x"E000B8",
   x"3C013B", x"010238", x"B0009E", x"01C082", x"100141",
   x"018000", x"100172", x"4000B4", x"100172", x"B00051",
   x"480000", x"B00030", x"B00059", x"000000", x"000000",
   x"000000", x"480001", x"B00051", x"B00030", x"B00059",
   x"000000", x"880002", x"000000", x"000000", x"B00051",
   x"01FFFC", x"C080B5", x"33011D", x"010230", x"B0009E",
   x"01C082", x"100141", x"010001", x"B0009E", x"013080",
   x"100141", x"010001", x"C08133", x"B0003F", x"280000",
   x"010001", x"C08135", x"010010", x"50812C", x"B0003F",
   x"280000", x"B00030", x"B00053", x"B0005B", x"000000",
   x"000000", x"000000", x"000000", x"B00053", x"40009E",
   x"B00030", x"B00051", x"B00059", x"000000", x"000000",
   x"000000", x"000000", x"B00051", x"B00040", x"280000",
   x"B00030", x"B00053", x"B0005B", x"000000", x"000000",
   x"000000", x"000000", x"B00053", x"B00041", x"B00045",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"400030", x"B0009F", x"000000",
   x"B00041", x"280000", x"400041", x"400045", x"000000",
   x"000000", x"000000", x"000000", x"400041", x"280000",
   x"B00030", x"B00051", x"B00059", x"000000", x"000000",
   x"000000", x"000000", x"B00051", x"280000", x"4000A5",
   x"B80000", x"4000A6", x"B80001", x"4000A7", x"B80002",
   x"4000A2", x"B80003", x"4000A3", x"B80004", x"4000A4",
   x"B80005", x"4000B6", x"B80006", x"280000", x"490003",
   x"B80000", x"490004", x"B80001", x"490005", x"B80002",
   x"4000A2", x"B80003", x"4000A3", x"B80004", x"4000A4",
   x"B80005", x"4000B6", x"B80006", x"280000", x"010001",
   x"060000", x"B80007", x"010800", x"060000", x"B80008",
   x"010604", x"060000", x"B80009", x"010002", x"060000",
   x"B8000A", x"4000A2", x"B8000B", x"4000A3", x"B8000C",
   x"4000A4", x"B8000D", x"4000A8", x"B8000E", x"4000A9",
   x"B8000F", x"49000B", x"B80010", x"49000C", x"B80011",
   x"49000D", x"B80012", x"49000E", x"B80013", x"49000F",
   x"B80014", x"280000", x"014500", x"060000", x"B80007",
   x"010000", x"060000", x"B80008", x"010000", x"060000",
   x"B80009", x"014000", x"060000", x"B8000A", x"014011",
   x"060000", x"B8000B", x"010000", x"060000", x"B8000C",
   x"4000A8", x"B8000D", x"4000AA", x"B8000E", x"4000AA",
   x"B8000F", x"4000AB", x"B80010", x"280000", x"014500",
   x"060000", x"B80007", x"010000", x"060000", x"B80008",
   x"010000", x"060000", x"B80009", x"014000", x"060000",
   x"B8000A", x"014011", x"060000", x"B8000B", x"010000",
   x"060000", x"B8000C", x"49000D", x"B8000F", x"49000E",
   x"B80010", x"4000A8", x"B8000D", x"4000A9", x"B8000E",
   x"280000", x"010000", x"060000", x"B80011", x"010000",
   x"060000", x"B80012", x"280000", x"490011", x"B80012",
   x"4000D8", x"B80011", x"010000", x"060000", x"B80014",
   x"280000", x"010044", x"060000", x"B80011", x"010043",
   x"060000", x"B80012", x"010134", x"060000", x"B80013",
   x"010000", x"060000", x"B80014", x"280000", x"010101",
   x"060000", x"B80015", x"010600", x"060000", x"B80016",
   x"4000BC", x"B80017", x"4000BD", x"B80018", x"010001",
   x"060000", x"B80019", x"018000", x"060000", x"B8001A",
   x"4000A8", x"B8001B", x"4000A9", x"B8001C", x"010000",
   x"060000", x"B8001D", x"010000", x"060000", x"B8001E",
   x"4000AA", x"B8001F", x"4000AB", x"B80020", x"010000",
   x"060000", x"B80021", x"010000", x"060000", x"B80022",
   x"4000A2", x"B80023", x"4000A3", x"B80024", x"4000A4",
   x"B80025", x"280000", x"1003E9", x"015A00", x"B00154",
   x"015A01", x"B0015C", x"015A02", x"B0011C", x"015A03",
   x"B00100", x"015A04", x"B00165", x"015A06", x"B00124",
   x"015A07", x"B0013C", x"016F48", x"B00158", x"017473",
   x"B00159", x"016F4D", x"B0015A", x"013274", x"B0015B",
   x"01534B", x"B00160", x"01385A", x"B00161", x"013538",
   x"B00162", x"010031", x"B00163", x"017445", x"B00120",
   x"016568", x"B00121", x"014572", x"B00122", x"015045",
   x"B00123", x"015046", x"B00104", x"014147", x"B00105",
   x"016C46", x"B00106", x"016873", x"B00107", x"016954",
   x"B00169", x"01656D", x"B0016A", x"017372", x"B0016B",
   x"010000", x"B0016C", x"01424C", x"B00128", x"013150",
   x"B00129", x"015236", x"B0012A", x"010057", x"B0012B",
   x"01424C", x"B00140", x"013150", x"B00141", x"015236",
   x"B00142", x"01004F", x"B00143", x"010130", x"870000",
   x"010008", x"B00137", x"010003", x"B0014C", x"01000F",
   x"B0014D", x"010001", x"B00081", x"010002", x"B00082",
   x"010003", x"B00083", x"010004", x"B00084", x"010005",
   x"B00085", x"010006", x"B00086", x"010007", x"B00087",
   x"010008", x"B00088", x"010010", x"B0008A", x"01000F",
   x"B00091", x"018104", x"B00155", x"010010", x"B00156",
   x"018102", x"B0015D", x"010008", x"B0015E", x"018E02",
   x"B0011D", x"010007", x"B0011E", x"018F04", x"B00101",
   x"018200", x"B00102", x"018202", x"B00166", x"010004",
   x"B00167", x"018202", x"B00125", x"010004", x"B00126",
   x"010202", x"B0013D", x"010004", x"B0013E", x"0100FF",
   x"B0008C", x"01FF00", x"B0008D", x"01FFFC", x"B0008E",
   x"010100", x"B0008F", x"011100", x"B00090", x"010400",
   x"B00092", x"010800", x"B00093", x"010C00", x"B00094",
   x"011000", x"B00095", x"011800", x"B00097", x"011C00",
   x"B00098", x"010100", x"B00099", x"010200", x"B0009A",
   x"01000F", x"B000EA", x"010060", x"060000", x"B000A2",
   x"011B10", x"060000", x"B000A3", x"010000", x"060000",
   x"B000A4", x"01FF00", x"060000", x"B000A5", x"010000",
   x"060000", x"B000A6", x"010000", x"060000", x"B000A7",
   x"016A2D", x"060000", x"B000D8", x"010044", x"060000",
   x"B000DA", x"010600", x"B000B9", x"010600", x"B000B8",
   x"0104B1", x"B000BB", x"0107FB", x"B000BA", x"01FFFF",
   x"B0007D", x"280000", x"010003", x"70003F", x"B0014E",
   x"E00081", x"3202FF", x"E00081", x"32030C", x"000000",
   x"000000", x"20035A", x"010011", x"B000D5", x"1007C8",
   x"4000D4", x"060000", x"B000A8", x"010010", x"B000D5",
   x"1007C8", x"4000D4", x"060000", x"B000A9", x"200360",
   x"1003FB", x"4000D0", x"B000BC", x"4000D1", x"B000BD",
   x"0104B6", x"840000", x"010148", x"B000B4", x"1003D9",
   x"010800", x"060000", x"B000B6", x"01FFFF", x"B000AA",
   x"B000AB", x"B000A5", x"B000A6", x"B000A7", x"010000",
   x"B000A8", x"B000A9", x"014011", x"060000", x"B8000B",
   x"10017B", x"1001BA", x"4000B4", x"060000", x"B80008",
   x"01000E", x"C080B4", x"1001FF", x"10020C", x"10010D",
   x"0103E8", x"B0009D", x"010001", x"100410", x"01FFFF",
   x"C0809D", x"32030C", x"4000AC", x"33033A", x"400031",
   x"330331", x"000000", x"000000", x"01017F", x"850000",
   x"10009E", x"320331", x"010180", x"850000", x"000000",
   x"000000", x"010800", x"060000", x"E90006", x"330331",
   x"49000B", x"E00090", x"70008D", x"330331", x"490012",
   x"E000DA", x"330331", x"490017", x"E000BC", x"330331",
   x"490018", x"E000BD", x"330331", x"49001D", x"B000A8",
   x"49001E", x"B000A9", x"200360", x"01C0A8", x"060000",
   x"B000A8", x"010179", x"060000", x"B000A9", x"280000",
   x"000000", x"010000", x"B00032", x"01000A", x"100410",
   x"010001", x"B00032", x"01000A", x"100410", x"010001",
   x"B0009E", x"01C026", x"100141", x"01000A", x"100410",
   x"010000", x"B0009E", x"01C026", x"100141", x"01000A",
   x"100410", x"013014", x"100154", x"40009F", x"060000",
   x"B000A2", x"01C012", x"100154", x"40009F", x"060000",
   x"B000A3", x"013010", x"100154", x"40009F", x"060000",
   x"B000A4", x"014000", x"B0009E", x"013084", x"100141",
   x"0101EE", x"B0009E", x"013070", x"100141", x"014000",
   x"B0009E", x"01C086", x"100141", x"010001", x"B0009E",
   x"01309C", x"100141", x"017CE0", x"B0009E", x"013074",
   x"100141", x"010016", x"B0009E", x"01C076", x"100141",
   x"010230", x"B0009E", x"01C082", x"100141", x"0120FF",
   x"B0009E", x"01C0F6", x"100141", x"01FFFF", x"B0009E",
   x"01C092", x"100141", x"012800", x"B0009E", x"013090",
   x"100141", x"0101EF", x"B0009E", x"013070", x"100141",
   x"017CE1", x"B0009E", x"013074", x"100141", x"4000A4",
   x"B000CC", x"B000CD", x"4000A3", x"B000CE", x"B000CF",
   x"000000", x"000000", x"000000", x"280000", x"010008",
   x"B000D5", x"010000", x"860000", x"1007C8", x"4000D4",
   x"BA0144", x"010001", x"C080D5", x"820000", x"E00087",
   x"3C03CE", x"8A0001", x"000000", x"2003C3", x"010014",
   x"B000D5", x"1007C8", x"4000D4", x"B00136", x"B0007B",
   x"100899", x"010004", x"C000E6", x"508102", x"280000",
   x"0B0000", x"B0009C", x"0104B6", x"860000", x"010000",
   x"BA0000", x"000000", x"000000", x"000000", x"01FFFF",
   x"8A0001", x"C0809C", x"3303DD", x"000000", x"000000",
   x"280000", x"010080", x"860000", x"010000", x"BA0000",
   x"000000", x"000000", x"000000", x"8A0001", x"820000",
   x"040000", x"040000", x"040000", x"040000", x"040000",
   x"3C03EB", x"000000", x"000000", x"280000", x"019069",
   x"A000CC", x"C000CD", x"B000CC", x"080000", x"D00080",
   x"B000CD", x"014650", x"A000CE", x"C000CF", x"B000CE",
   x"080000", x"D00080", x"B000CF", x"4000CE", x"B000D0",
   x"000000", x"4000CF", x"C000CD", x"B000D1", x"280000",
   x"B000BE", x"0137CE", x"B000BF", x"000000", x"000000",
   x"01FFFF", x"C080BF", x"000000", x"000000", x"330415",
   x"01FFFF", x"C080BE", x"330411", x"000000", x"000000",
   x"280000", x"011100", x"B00068", x"01FFFF", x"B00060",
   x"B00061", x"B0006D", x"000000", x"000000", x"000000",
   x"011104", x"B00068", x"01FFFF", x"B00060", x"B00061",
   x"B0006D", x"000000", x"000000", x"000000", x"011108",
   x"B00068", x"01FFFF", x"B00060", x"B00061", x"B0006D",
   x"000000", x"000000", x"000000", x"01110C", x"B00068",
   x"01FFFF", x"B00060", x"B00061", x"B0006D", x"000000",
   x"000000", x"000000", x"011000", x"B00068", x"010000",
   x"B00060", x"B00061", x"B0006D", x"000000", x"000000",
   x"000000", x"011004", x"B00068", x"010000", x"B00060",
   x"B00061", x"B0006D", x"000000", x"000000", x"000000",
   x"011008", x"B00068", x"010000", x"B00060", x"B00061",
   x"B0006D", x"000000", x"000000", x"000000", x"01100C",
   x"B00068", x"010000", x"B00060", x"B00061", x"B0006D",
   x"000000", x"000000", x"000000", x"280000", x"810000",
   x"C000DC", x"B000DD", x"800000", x"B000DE", x"490000",
   x"B000DF", x"000000", x"890001", x"01007F", x"7000DF",
   x"3204B6", x"B0009B", x"013C00", x"7000DF", x"3304D1",
   x"010300", x"7000DF", x"E0009A", x"3304B6", x"014000",
   x"7000DF", x"320484", x"490000", x"B00157", x"890001",
   x"200485", x"400157", x"B00068", x"018000", x"7000DF",
   x"33049A", x"B0006C", x"800000", x"E000BA", x"3C04BE",
   x"4000DF", x"B0006E", x"400060", x"B80000", x"400061",
   x"B80001", x"01FFFF", x"C0809B", x"880002", x"330489",
   x"400068", x"B00157", x"2004AB", x"490000", x"B00060",
   x"490001", x"B00061", x"810000", x"E000BB", x"3C04BE",
   x"B0006D", x"890002", x"4000DF", x"B0006E", x"01FFFF",
   x"C0809B", x"33049A", x"000000", x"400068", x"B00157",
   x"810000", x"E000DD", x"38046E", x"010001", x"C08131",
   x"010000", x"B00139", x"800000", x"E000DE", x"040000",
   x"20007B", x"010001", x"50812C", x"01FFFF", x"E0012D",
   x"3204CD", x"010001", x"C0812D", x"2004CD", x"010002",
   x"50812C", x"01FFFF", x"E0012E", x"3204CD", x"010001",
   x"C0812E", x"2004CD", x"010004", x"50812C", x"01FFFF",
   x"E0012F", x"3204CD", x"010001", x"C0812F", x"010000",
   x"B00139", x"8F0000", x"20007B", x"011C00", x"7000DF",
   x"E00095", x"3205A1", x"011C00", x"7000DF", x"E00092",
   x"320666", x"011C00", x"7000DF", x"E00093", x"3206C3",
   x"011C00", x"7000DF", x"E00094", x"32071E", x"011C00",
   x"7000DF", x"E00098", x"3204EF", x"011C00", x"7000DF",
   x"E00097", x"320529", x"011C00", x"7000DF", x"320653",
   x"000000", x"000000", x"2004B6", x"012000", x"7000DF",
   x"330516", x"010300", x"7000DF", x"E00099", x"3304B6",
   x"014000", x"7000DF", x"3204FD", x"490000", x"B0013F",
   x"890001", x"2004FF", x"000000", x"40013F", x"0B0000",
   x"860000", x"018000", x"7000DF", x"3304C6", x"820000",
   x"E0008A", x"3C04BE", x"4A0144", x"B80000", x"010080",
   x"7000DF", x"32050F", x"010002", x"C0813F", x"8A0001",
   x"01FFFF", x"C0809B", x"880001", x"330504", x"000000",
   x"000000", x"2004AB", x"100797", x"820000", x"E00088",
   x"3C04BE", x"4A013C", x"B80000", x"010080", x"7000DF",
   x"320522", x"010002", x"C080E2", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"330517", x"000000", x"000000",
   x"2004AB", x"012000", x"7000DF", x"33058E", x"010300",
   x"7000DF", x"E00099", x"3304B6", x"014000", x"7000DF",
   x"320537", x"490000", x"B00127", x"890001", x"200538",
   x"400127", x"0B0000", x"860000", x"018000", x"7000DF",
   x"330565", x"820000", x"E0008A", x"3C04BE", x"820000",
   x"E000EA", x"330556", x"010001", x"B00022", x"000000",
   x"000000", x"010001", x"B00021", x"000000", x"000000",
   x"000000", x"010000", x"B00021", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"400020", x"B80000",
   x"200558", x"4A012C", x"B80000", x"010080", x"7000DF",
   x"32055E", x"010002", x"C08127", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"33053D", x"000000", x"000000",
   x"2004AB", x"820000", x"E0008A", x"3C04BE", x"820000",
   x"E000EA", x"330578", x"010000", x"B00022", x"490000",
   x"B00020", x"000000", x"000000", x"010001", x"B00021",
   x"000000", x"000000", x"010000", x"B00021", x"20057A",
   x"490000", x"BA012C", x"010080", x"7000DF", x"320580",
   x"010002", x"C08127", x"8A0001", x"01FFFF", x"C0809B",
   x"890001", x"330565", x"400136", x"B0007B", x"01012C",
   x"B000A0", x"01001F", x"700137", x"0B0000", x"C000A0",
   x"870000", x"2004AB", x"100797", x"820000", x"E00088",
   x"3C04BE", x"4A0124", x"B80000", x"010080", x"7000DF",
   x"32059A", x"010002", x"C080E2", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"33058F", x"000000", x"000000",
   x"2004AB", x"012000", x"7000DF", x"330640", x"010300",
   x"7000DF", x"E00099", x"3304B6", x"014000", x"7000DF",
   x"3205AF", x"490000", x"B00168", x"890001", x"2005B0",
   x"400168", x"0B0000", x"860000", x"018000", x"7000DF",
   x"3305FC", x"820000", x"E0008A", x"3C04BE", x"820000",
   x"E00088", x"3805BE", x"4A016E", x"000000", x"2005EE",
   x"820000", x"3305C3", x"40007C", x"000000", x"2005EE",
   x"820000", x"E00081", x"3305C9", x"40016F", x"000000",
   x"2005EE", x"820000", x"E00082", x"3305CF", x"4A016E",
   x"000000", x"2005EE", x"820000", x"E00083", x"3305D6",
   x"010001", x"B000C1", x"1007A9", x"2005EE", x"820000",
   x"E00084", x"3305DD", x"010002", x"B000C1", x"1007A9",
   x"2005EE", x"820000", x"E00085", x"3305E4", x"010004",
   x"B000C1", x"1007A9", x"2005EE", x"820000", x"E00086",
   x"3305EB", x"010008", x"B000C1", x"1007A9", x"2005EE",
   x"010010", x"B000C1", x"1007A9", x"B80000", x"010080",
   x"7000DF", x"3205F5", x"010002", x"C08168", x"8A0001",
   x"01FFFF", x"C0809B", x"880001", x"3305B5", x"000000",
   x"000000", x"2004AB", x"820000", x"E0008A", x"3C04BE",
   x"490000", x"BA016E", x"820000", x"330606", x"000000",
   x"000000", x"200633", x"820000", x"E00081", x"33060E",
   x"40007C", x"B000C6", x"000000", x"1007C1", x"200633",
   x"820000", x"E00082", x"330614", x"000000", x"000000",
   x"200633", x"820000", x"E00083", x"33061B", x"010001",
   x"B000C1", x"1007A9", x"200633", x"820000", x"E00084",
   x"330622", x"010002", x"B000C1", x"1007A9", x"200633",
   x"820000", x"E00085", x"330629", x"010004", x"B000C1",
   x"1007A9", x"200633", x"820000", x"E00086", x"330630",
   x"010008", x"B000C1", x"1007A9", x"200633", x"010010",
   x"B000C1", x"1007A9", x"8A0001", x"010080", x"7000DF",
   x"320639", x"010002", x"C08168", x"01FFFF", x"C0809B",
   x"890001", x"3305FC", x"000000", x"000000", x"2004AB",
   x"100797", x"820000", x"E00088", x"3C04BE", x"4A0165",
   x"B80000", x"010080", x"7000DF", x"32064C", x"010002",
   x"C080E2", x"8A0001", x"01FFFF", x"C0809B", x"880001",
   x"330641", x"000000", x"000000", x"2004AB", x"100797",
   x"820000", x"E00088", x"3C04BE", x"4A0154", x"B80000",
   x"010080", x"7000DF", x"32065F", x"010002", x"C080E2",
   x"8A0001", x"01FFFF", x"C0809B", x"880001", x"330654",
   x"000000", x"000000", x"2004AB", x"012000", x"7000DF",
   x"3306B0", x"010300", x"7000DF", x"E00099", x"3304B6",
   x"014000", x"7000DF", x"320674", x"490000", x"B0015F",
   x"890001", x"200675", x"40015F", x"0B0000", x"860000",
   x"010002", x"70015F", x"32067E", x"01C000", x"50015F",
   x"B000E0", x"200681", x"013000", x"50015F", x"B000E0",
   x"018000", x"7000DF", x"33069A", x"010F00", x"7000E0",
   x"3304BE", x"000000", x"4000E0", x"100154", x"40009F",
   x"B80000", x"010080", x"7000DF", x"320693", x"010002",
   x"C0815F", x"010002", x"C080E0", x"01FFFF", x"C0809B",
   x"880001", x"330684", x"000000", x"000000", x"2004AB",
   x"010F00", x"7000E0", x"3304BE", x"490000", x"B0009E",
   x"4000E0", x"100141", x"010080", x"7000DF", x"3206A9",
   x"010002", x"C0815F", x"010002", x"C080E0", x"8A0001",
   x"01FFFF", x"C0809B", x"890001", x"33069A", x"000000",
   x"000000", x"2004AB", x"100797", x"820000", x"E00088",
   x"3C04BE", x"4A015C", x"B80000", x"010080", x"7000DF",
   x"3206BC", x"010002", x"C080E2", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"3306B1", x"000000", x"000000",
   x"2004AB", x"012000", x"7000DF", x"33070B", x"010300",
   x"7000DF", x"E00099", x"3304B6", x"014000", x"7000DF",
   x"3206D1", x"490000", x"B0011F", x"890001", x"2006D2",
   x"40011F", x"0B0000", x"860000", x"B000D5", x"018000",
   x"7000DF", x"3306EE", x"01FFC0", x"7000D5", x"3304BE",
   x"000000", x"000000", x"1007C8", x"4000D4", x"B80000",
   x"010080", x"7000DF", x"3206E7", x"010002", x"C0811F",
   x"010001", x"C080D5", x"01FFFF", x"C0809B", x"880001",
   x"3306D8", x"000000", x"000000", x"2004AB", x"013602",
   x"E00139", x"3206F7", x"015A02", x"E00139", x"3304C6",
   x"01000F", x"E000D5", x"3C04C6", x"01FFC0", x"7000D5",
   x"3304BE", x"490000", x"B000D3", x"1007D1", x"010080",
   x"7000DF", x"320704", x"010002", x"C0811F", x"010001",
   x"C080D5", x"01FFFF", x"C0809B", x"890001", x"3306EE",
   x"000000", x"000000", x"2004AB", x"100797", x"820000",
   x"E00088", x"3C04BE", x"4A011C", x"B80000", x"010080",
   x"7000DF", x"320717", x"010002", x"C080E2", x"8A0001",
   x"01FFFF", x"C0809B", x"880001", x"33070C", x"000000",
   x"000000", x"2004AB", x"012000", x"7000DF", x"330784",
   x"014000", x"7000DF", x"320728", x"490000", x"B00103",
   x"890001", x"200729", x"400103", x"860000", x"012000",
   x"7000DF", x"330784", x"010300", x"7000DF", x"E0009A",
   x"3304B6", x"018000", x"7000DF", x"33075A", x"800000",
   x"E000BA", x"3C04BE", x"400103", x"320740", x"E00084",
   x"320746", x"E00084", x"32074C", x"000000", x"000000",
   x"2004BE", x"1008C7", x"4000E4", x"B80000", x"4000E5",
   x"B80001", x"200752", x"100880", x"010004", x"C080E4",
   x"010000", x"D080E5", x"20074E", x"1008C7", x"100899",
   x"4000E6", x"B80000", x"4000E7", x"B80001", x"01FFFF",
   x"C0809B", x"000000", x"880002", x"330734", x"000000",
   x"000000", x"2004AB", x"400103", x"320763", x"E00084",
   x"320771", x"E00088", x"320769", x"000000", x"000000",
   x"2004BE", x"1008C7", x"490000", x"B000E4", x"490001",
   x"B000E5", x"20077D", x"1008C7", x"015A03", x"E00139",
   x"3304C6", x"000000", x"000000", x"1008BC", x"20077D",
   x"015A03", x"E00139", x"3304C6", x"490000", x"B000E6",
   x"490001", x"B000E7", x"1008A6", x"010004", x"C080E4",
   x"010000", x"D080E5", x"01FFFF", x"C0809B", x"890002",
   x"33075A", x"000000", x"000000", x"2004AB", x"100797",
   x"820000", x"E00088", x"3C04BE", x"4A0100", x"B80000",
   x"010080", x"7000DF", x"320790", x"010003", x"C080E2",
   x"8A0001", x"01FFFF", x"C0809B", x"880001", x"330785",
   x"000000", x"000000", x"2004AB", x"010300", x"7000DF",
   x"E00099", x"3304B6", x"018000", x"7000DF", x"3304C6",
   x"014000", x"7000DF", x"3207A5", x"490000", x"B000E2",
   x"890001", x"2007A6", x"4000E2", x"0B0000", x"860000",
   x"280000", x"010000", x"B000C5", x"40007C", x"B000C4",
   x"400070", x"7000C1", x"B000C3", x"400070", x"7000C1",
   x"B000C2", x"3207B6", x"4000C3", x"3207BF", x"4000C2",
   x"B000C3", x"40007C", x"E000C4", x"B000C5", x"E00170",
   x"3807B0", x"010020", x"50812C", x"4000C5", x"280000",
   x"40007C", x"E000C6", x"E0016F", x"3807C1", x"000000",
   x"000000", x"280000", x"100842", x"010006", x"100812",
   x"4000D5", x"100825", x"10084D", x"B000D4", x"100849",
   x"280000", x"100842", x"010004", x"100812", x"01003F",
   x"100825", x"100849", x"100842", x"010005", x"100812",
   x"4000D5", x"100825", x"1007FE", x"100804", x"4000D3",
   x"10085E", x"100849", x"100871", x"100842", x"010004",
   x"100812", x"010000", x"100825", x"100849", x"280000",
   x"010002", x"5080D2", x"280000", x"01FFFD", x"7080D2",
   x"280000", x"010001", x"5080D2", x"280000", x"01FFFE",
   x"7080D2", x"280000", x"3307FB", x"000000", x"000000",
   x"01FFFB", x"7080D2", x"280000", x"010004", x"5080D2",
   x"280000", x"010020", x"5080D2", x"280000", x"01FFDF",
   x"7080D2", x"280000", x"B0009E", x"01C022", x"100141",
   x"280000", x"01C022", x"100154", x"010008", x"70009F",
   x"280000", x"1007E9", x"100804", x"1007EC", x"100804",
   x"280000", x"B000A0", x"000000", x"000000", x"010004",
   x"7000A0", x"1007F5", x"100804", x"10080D", x"010002",
   x"7000A0", x"1007F5", x"100804", x"10080D", x"010001",
   x"7000A0", x"1007F5", x"100804", x"10080D", x"280000",
   x"B000A0", x"010020", x"B000D6", x"000000", x"000000",
   x"4000A0", x"7000D6", x"1007F5", x"100804", x"4000D6",
   x"C00080", x"050000", x"B000D6", x"1007E9", x"100804",
   x"1007EC", x"4000D6", x"33083B", x"000000", x"000000",
   x"100801", x"20083C", x"1007FE", x"100804", x"4000D6",
   x"33082A", x"000000", x"000000", x"280000", x"010000",
   x"B000D2", x"100804", x"010031", x"B000D2", x"100804",
   x"280000", x"010000", x"B000D2", x"100804", x"280000",
   x"B000A0", x"018000", x"B000D6", x"10080D", x"100808",
   x"320855", x"4000D6", x"5080A0", x"10080D", x"4000D6",
   x"C00080", x"050000", x"B000D6", x"330851", x"4000A0",
   x"000000", x"280000", x"B000A0", x"018000", x"B000D6",
   x"000000", x"000000", x"4000A0", x"7000D6", x"1007F5",
   x"100804", x"10080D", x"4000D6", x"C00080", x"050000",
   x"B000D6", x"000000", x"330863", x"000000", x"000000",
   x"280000", x"01C350", x"B000A0", x"010011", x"B000D2",
   x"100804", x"100808", x"33087E", x"01FFFF", x"C080A0",
   x"330876", x"000000", x"000000", x"2004C6", x"100849",
   x"280000", x"01AA02", x"E000E8", x"32088A", x"01AA02",
   x"B000E8", x"010000", x"B0007D", x"010003", x"1008E5",
   x"1008EE", x"010000", x"1008E5", x"B000E6", x"010000",
   x"1008E5", x"060000", x"5080E6", x"010000", x"1008E5",
   x"B000E7", x"010000", x"1008E5", x"060000", x"5080E7",
   x"280000", x"010000", x"B0007D", x"0100AB", x"1008E5",
   x"1008EE", x"010000", x"1008E5", x"B000E6", x"010000",
   x"B000E7", x"01FFFF", x"B0007D", x"280000", x"01AA03",
   x"E000E8", x"3208B1", x"01AA03", x"B000E8", x"100900",
   x"010000", x"B0007D", x"010002", x"1008E5", x"1008EE",
   x"4000E6", x"1008E5", x"4000E6", x"060000", x"1008E5",
   x"4000E7", x"1008E5", x"4000E7", x"060000", x"1008E5",
   x"280000", x"100900", x"010000", x"B0007D", x"0100D8",
   x"1008E5", x"1008EE", x"010BB8", x"1008D4", x"01AA01",
   x"B000E8", x"280000", x"01AA03", x"E000E8", x"3208CF",
   x"01FFFF", x"B0007D", x"01AA01", x"B000E8", x"280000",
   x"010005", x"1008D4", x"01AA01", x"B000E8", x"280000",
   x"B0009C", x"01FFFF", x"B0007D", x"1008F6", x"700081",
   x"3208E3", x"000000", x"010001", x"100410", x"01FFFF",
   x"C0809C", x"3308D7", x"000000", x"000000", x"2004C6",
   x"100907", x"280000", x"B0007E", x"000000", x"010002",
   x"70007D", x"3308E6", x"0100FF", x"70007E", x"B000E9",
   x"280000", x"4000E5", x"1008E5", x"4000E4", x"060000",
   x"1008E5", x"4000E4", x"1008E5", x"280000", x"010000",
   x"B0007D", x"010005", x"1008E5", x"010000", x"1008E5",
   x"01FFFF", x"B0007D", x"4000E9", x"280000", x"010000",
   x"B0007D", x"010006", x"1008E5", x"010001", x"B0007D",
   x"280000", x"010000", x"B0007D", x"010004", x"1008E5",
   x"010001", x"B0007D", x"280000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"00ABCD");

signal daddr: std_logic_vector(11 downto 0);

begin
   aetherhm2: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (we = '1') then
            RAM(conv_integer(addr)) <= din;
         end if;
         daddr <= addr;
      end if; -- clk 
   end process;

   dout <= RAM(conv_integer(daddr));
end;
