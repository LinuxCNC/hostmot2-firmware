library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from sslbp.bin
-- On 11/ 8/2010

entity sslbp is
	port (
	addra: in std_logic_vector(10 downto 0);
	addrb: in std_logic_vector(10 downto 0);
	clk: in std_logic;
	dina: in std_logic_vector(15 downto 0);
	douta: out std_logic_vector(15 downto 0);
	doutb: out std_logic_vector(15 downto 0);
	wea: in std_logic);
end sslbp;

architecture syn of sslbp is
   type ram_type is array (0 to 2047) of std_logic_vector(15 downto 0);
   signal RAM : ram_type := 
   (
   x"0000", x"0000", x"0100", x"B028", x"B054", x"B049", x"B04C", x"0101",
   x"B029", x"01FF", x"B02A", x"0155", x"B02B", x"01AA", x"B402", x"7434",
   x"B04A", x"0138", x"B008", x"0149", x"B009", x"0132", x"B00A", x"0130",
   x"B00B", x"0137", x"B00C", x"0149", x"B00D", x"0136", x"B00E", x"0134",
   x"B00F", x"0112", x"B000", x"0101", x"B002", x"010B", x"B003", x"0108",
   x"B001", x"01D8", x"B006", x"704A", x"B007", x"0180", x"0800", x"0100",
   x"0A00", x"0002", x"704A", x"B045", x"01A0", x"B818", x"0125", x"B819",
   x"0126", x"B81A", x"0100", x"B81B", x"0C20", x"7045", x"E029", x"B045",
   x"2034", x"0100", x"B049", x"0100", x"B04C", x"B400", x"7049", x"3563",
   x"0180", x"0800", x"0100", x"0A00", x"0180", x"0880", x"0101", x"0A80",
   x"0180", x"0900", x"0104", x"0B00", x"0100", x"0980", x"0106", x"0B80",
   x"0101", x"B052", x"01FE", x"B053", x"704A", x"B044", x"0180", x"A801",
   x"2526", x"7054", x"A052", x"3526", x"016B", x"C800", x"0E80", x"0000",
   x"0000", x"0000", x"1800", x"11B6", x"11BB", x"11BF", x"11CD", x"11D5",
   x"11E0", x"1513", x"151D", x"1216", x"1220", x"1227", x"122F", x"1236",
   x"123B", x"1243", x"124A", x"1255", x"125D", x"1264", x"126E", x"1275",
   x"127F", x"1286", x"1290", x"1297", x"12C3", x"1309", x"1319", x"1320",
   x"132C", x"1333", x"133C", x"134C", x"1353", x"138F", x"139F", x"13A6",
   x"13B6", x"13BD", x"13C9", x"13D0", x"13D9", x"13E5", x"13EC", x"142B",
   x"143B", x"10F1", x"10FB", x"1102", x"10AB", x"10C0", x"10CE", x"12EF",
   x"12FF", x"118C", x"119C", x"1145", x"115A", x"1168", x"1446", x"14B5",
   x"14C3", x"1524", x"1525", x"7057", x"A052", x"30BF", x"0003", x"0003",
   x"678B", x"705C", x"67C0", x"79A0", x"67C0", x"79A1", x"67C0", x"79A2",
   x"67C0", x"79A3", x"67C0", x"67C3", x"66A0", x"0132", x"B800", x"1526",
   x"6759", x"50C4", x"0131", x"B800", x"0108", x"6705", x"30CD", x"40CB",
   x"0131", x"B800", x"10CD", x"0133", x"B800", x"1526", x"7880", x"B9C0",
   x"7881", x"B9C1", x"7882", x"B9C2", x"7883", x"B9C3", x"8882", x"30DB",
   x"0101", x"8802", x"B802", x"7886", x"B9A0", x"7887", x"B9A1", x"7884",
   x"B9A2", x"7885", x"B9A3", x"7057", x"A053", x"B057", x"7802", x"20EE",
   x"7058", x"A053", x"B058", x"7059", x"A053", x"B059", x"0131", x"B800",
   x"1526", x"0101", x"B809", x"678B", x"01DF", x"67C0", x"67C3", x"012F",
   x"B800", x"66A0", x"1526", x"6759", x"0101", x"6705", x"3101", x"0130",
   x"B800", x"1526", x"015A", x"E880", x"2117", x"017F", x"A802", x"B802",
   x"7055", x"A053", x"B055", x"7056", x"A053", x"B056", x"7057", x"A052",
   x"3114", x"0131", x"B800", x"1116", x"012E", x"B800", x"1144", x"0101",
   x"C804", x"511D", x"B804", x"0003", x"1132", x"7809", x"E804", x"4132",
   x"0180", x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801",
   x"312C", x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940",
   x"0100", x"B950", x"0102", x"8801", x"B801", x"7059", x"A053", x"B059",
   x"0180", x"A801", x"313E", x"7056", x"A053", x"B056", x"0120", x"8802",
   x"B802", x"B940", x"0100", x"B950", x"1526", x"7057", x"A052", x"3159",
   x"0003", x"0003", x"678B", x"705C", x"67C0", x"79A0", x"67C0", x"79A1",
   x"67C0", x"79A2", x"67C0", x"0100", x"67C0", x"67C3", x"66A0", x"0139",
   x"B800", x"1526", x"6759", x"515E", x"0138", x"B800", x"0108", x"6705",
   x"3167", x"4165", x"0138", x"B800", x"1167", x"013A", x"B800", x"1526",
   x"7880", x"B9A0", x"7881", x"B9A1", x"7882", x"B9A2", x"0108", x"A883",
   x"3174", x"0101", x"8802", x"B802", x"0100", x"B9A3", x"7884", x"B9C0",
   x"7885", x"B9C1", x"7886", x"B9C2", x"7887", x"B9C3", x"7057", x"A053",
   x"B057", x"7802", x"2189", x"7058", x"A053", x"B058", x"7059", x"A053",
   x"B059", x"0138", x"B800", x"1526", x"678B", x"705C", x"67C0", x"0100",
   x"67C0", x"0100", x"67C0", x"0100", x"67C0", x"0100", x"67C0", x"67C3",
   x"0137", x"B800", x"66A0", x"1526", x"6759", x"0108", x"6705", x"31B5",
   x"017F", x"A802", x"B802", x"7055", x"A053", x"B055", x"7056", x"A053",
   x"B056", x"7057", x"A052", x"31AF", x"0138", x"B800", x"11B5", x"0128",
   x"B812", x"0100", x"B813", x"0136", x"B800", x"1526", x"66A5", x"B940",
   x"0101", x"B800", x"1526", x"66A0", x"0102", x"B800", x"1526", x"7422",
   x"E810", x"B031", x"7423", x"F811", x"B032", x"7812", x"E031", x"7813",
   x"F032", x"41CC", x"0103", x"B800", x"1526", x"678B", x"01DF", x"67C0",
   x"67C3", x"0104", x"B800", x"66A0", x"1526", x"6759", x"51DA", x"0101",
   x"B800", x"11DF", x"0101", x"6705", x"31DF", x"0105", x"B800", x"1526",
   x"015A", x"E880", x"21E6", x"0106", x"B800", x"1215", x"0101", x"C804",
   x"51EC", x"B804", x"0003", x"1201", x"7809", x"E804", x"4201", x"0180",
   x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"31FB",
   x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100",
   x"B950", x"0102", x"8801", x"B801", x"7059", x"A053", x"B059", x"0180",
   x"A801", x"320D", x"7056", x"A053", x"B056", x"0120", x"8802", x"B802",
   x"B940", x"0100", x"B950", x"0101", x"B800", x"1526", x"678B", x"01E1",
   x"67C0", x"0100", x"67C0", x"67C3", x"0109", x"B800", x"66A0", x"1526",
   x"6759", x"0100", x"6705", x"3226", x"010A", x"B800", x"1526", x"678B",
   x"01C1", x"67C0", x"67C3", x"010B", x"B800", x"66A0", x"1526", x"6759",
   x"0101", x"6705", x"3235", x"010C", x"B800", x"1526", x"7880", x"223A",
   x"010D", x"B800", x"1526", x"678B", x"01BC", x"67C0", x"67C3", x"010E",
   x"B800", x"66A0", x"1526", x"6759", x"0104", x"6705", x"3249", x"010F",
   x"B800", x"1526", x"7880", x"B9A0", x"7881", x"B9A1", x"7882", x"B9A2",
   x"7883", x"B9A3", x"0110", x"B800", x"1526", x"678B", x"01D0", x"67C0",
   x"67C3", x"0111", x"B800", x"66A0", x"1526", x"6759", x"0101", x"6705",
   x"3263", x"0112", x"B800", x"1526", x"7880", x"B814", x"678B", x"01D1",
   x"67C0", x"67C3", x"0113", x"B800", x"66A0", x"1526", x"6759", x"0101",
   x"6705", x"3274", x"0114", x"B800", x"1526", x"7880", x"B815", x"678B",
   x"01D2", x"67C0", x"67C3", x"0115", x"B800", x"66A0", x"1526", x"6759",
   x"0101", x"6705", x"3285", x"0116", x"B800", x"1526", x"7880", x"B816",
   x"678B", x"01D3", x"67C0", x"67C3", x"0117", x"B800", x"66A0", x"1526",
   x"6759", x"0101", x"6705", x"3296", x"0118", x"B800", x"1526", x"0119",
   x"B800", x"7880", x"B817", x"7008", x"E814", x"B030", x"7009", x"F815",
   x"8030", x"B030", x"700A", x"F816", x"8030", x"B030", x"700B", x"F817",
   x"8030", x"22C2", x"0180", x"B80C", x"0109", x"E048", x"22B4", x"01BF",
   x"A802", x"B802", x"011A", x"B800", x"010F", x"E048", x"22C2", x"013E",
   x"A802", x"B802", x"7055", x"A053", x"B055", x"7056", x"A053", x"B056",
   x"013B", x"B800", x"1526", x"013F", x"B800", x"7880", x"B817", x"700C",
   x"E814", x"B030", x"700D", x"F815", x"8030", x"B030", x"700E", x"F816",
   x"8030", x"B030", x"700F", x"F817", x"8030", x"22EE", x"0174", x"B80C",
   x"0109", x"E048", x"22E0", x"01BF", x"A802", x"B802", x"0134", x"B800",
   x"010F", x"E048", x"22EE", x"013E", x"A802", x"B802", x"7055", x"A053",
   x"B055", x"7056", x"A053", x"B056", x"013B", x"B800", x"1526", x"678B",
   x"705C", x"67C0", x"0100", x"67C0", x"0100", x"67C0", x"0100", x"67C0",
   x"0108", x"67C0", x"67C3", x"0135", x"B800", x"66A0", x"1526", x"6759",
   x"0108", x"6705", x"3308", x"01FE", x"A802", x"B802", x"0136", x"B800",
   x"1526", x"678B", x"0165", x"67C0", x"0154", x"67C0", x"0108", x"67C0",
   x"01FF", x"67C0", x"01FF", x"67C0", x"67C3", x"011B", x"B800", x"66A0",
   x"1526", x"6759", x"0100", x"6705", x"331F", x"011C", x"B800", x"1526",
   x"678B", x"0145", x"67C0", x"0154", x"67C0", x"0108", x"67C0", x"67C3",
   x"011D", x"B800", x"66A0", x"1526", x"6759", x"0102", x"6705", x"3332",
   x"011E", x"B800", x"1526", x"7880", x"8881", x"2339", x"011F", x"B800",
   x"133B", x"011C", x"B800", x"1526", x"7880", x"B05D", x"7881", x"B05E",
   x"678B", x"0145", x"67C0", x"0152", x"67C0", x"0108", x"67C0", x"67C3",
   x"0120", x"B800", x"66A0", x"1526", x"6759", x"0102", x"6705", x"3352",
   x"0121", x"B800", x"1526", x"0180", x"B9C0", x"0100", x"B9C1", x"7880",
   x"B9C2", x"7881", x"B9C3", x"7880", x"8881", x"2361", x"0122", x"B800",
   x"138E", x"0101", x"C808", x"5367", x"B808", x"0003", x"137C", x"7809",
   x"E808", x"437C", x"0180", x"8801", x"B801", x"7059", x"A053", x"B059",
   x"0180", x"A801", x"3376", x"7056", x"A053", x"B056", x"0120", x"8802",
   x"B802", x"B940", x"0100", x"B950", x"0140", x"8801", x"B801", x"7059",
   x"A053", x"B059", x"0180", x"A801", x"3388", x"7056", x"A053", x"B056",
   x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"1526", x"678B",
   x"0165", x"67C0", x"0160", x"67C0", x"0108", x"67C0", x"0100", x"67C0",
   x"0100", x"67C0", x"67C3", x"0123", x"B800", x"66A0", x"1526", x"6759",
   x"0100", x"6705", x"33A5", x"0124", x"B800", x"1526", x"678B", x"0165",
   x"67C0", x"0104", x"67C0", x"0108", x"67C0", x"01FF", x"67C0", x"01FF",
   x"67C0", x"67C3", x"0125", x"B800", x"66A0", x"1526", x"6759", x"0100",
   x"6705", x"33BC", x"0126", x"B800", x"1526", x"678B", x"0145", x"67C0",
   x"01FE", x"67C0", x"0108", x"67C0", x"67C3", x"0127", x"B800", x"66A0",
   x"1526", x"6759", x"0102", x"6705", x"33CF", x"0128", x"B800", x"1526",
   x"7880", x"8881", x"23D6", x"0126", x"B800", x"13D8", x"0129", x"B800",
   x"1526", x"678B", x"0145", x"67C0", x"0152", x"67C0", x"0108", x"67C0",
   x"67C3", x"012A", x"B800", x"66A0", x"1526", x"6759", x"0102", x"6705",
   x"33EB", x"012B", x"B800", x"1526", x"0180", x"B9C0", x"0100", x"B9C1",
   x"7880", x"B9C2", x"7881", x"B9C3", x"7880", x"8881", x"23FD", x"01FE",
   x"A802", x"B802", x"012C", x"B800", x"142A", x"0101", x"C808", x"5403",
   x"B808", x"0003", x"1418", x"7809", x"E808", x"4418", x"0180", x"8801",
   x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"3412", x"7056",
   x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950",
   x"0140", x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801",
   x"3424", x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940",
   x"0100", x"B950", x"1526", x"678B", x"0165", x"67C0", x"015C", x"67C0",
   x"0108", x"67C0", x"01F4", x"67C0", x"0101", x"67C0", x"67C3", x"012D",
   x"B800", x"66A0", x"1526", x"6759", x"0100", x"6705", x"3445", x"010F",
   x"B812", x"0100", x"B813", x"012E", x"B800", x"1526", x"7057", x"A052",
   x"34B4", x"0003", x"0003", x"678B", x"7980", x"B050", x"7981", x"B051",
   x"7983", x"B04F", x"67C0", x"0103", x"A04F", x"B046", x"C028", x"0101",
   x"B047", x"7046", x"3463", x"7047", x"0200", x"B047", x"7046", x"E029",
   x"B046", x"0001", x"1459", x"01BF", x"E04F", x"54A5", x"0104", x"A04F",
   x"346E", x"0003", x"7050", x"67C0", x"7051", x"67C0", x"0120", x"A04F",
   x"34A2", x"0100", x"B80A", x"0108", x"E047", x"2487", x"0003", x"79A0",
   x"67C0", x"79A1", x"67C0", x"79A2", x"67C0", x"79A3", x"67C0", x"79C0",
   x"67C0", x"79C1", x"67C0", x"79C2", x"67C0", x"79C3", x"67C0", x"0104",
   x"E047", x"2493", x"0003", x"79A0", x"67C0", x"79A1", x"67C0", x"79A2",
   x"67C0", x"79A3", x"67C0", x"0102", x"E047", x"249B", x"0003", x"79A0",
   x"67C0", x"79A1", x"67C0", x"0101", x"E047", x"24A1", x"0003", x"79A0",
   x"67C0", x"14A4", x"7047", x"B80A", x"14B0", x"0120", x"A04F", x"34AE",
   x"0003", x"79A0", x"67C0", x"0100", x"B80A", x"14B0", x"0101", x"B80A",
   x"67C3", x"66A0", x"013C", x"B800", x"1526", x"6759", x"54B9", x"013B",
   x"B800", x"780A", x"6705", x"34C2", x"44C0", x"013B", x"B800", x"14C2",
   x"013D", x"B800", x"1526", x"780A", x"B030", x"0001", x"0001", x"0108",
   x"E030", x"24DA", x"7880", x"B9A0", x"7881", x"B9A1", x"7882", x"B9A2",
   x"7883", x"B9A3", x"7884", x"B9C0", x"7885", x"B9C1", x"7886", x"B9C2",
   x"7887", x"B9C3", x"0104", x"E030", x"24EA", x"7880", x"B9A0", x"7881",
   x"B9A1", x"7882", x"B9A2", x"7883", x"B9A3", x"0100", x"B9C0", x"B9C1",
   x"B9C2", x"B9C3", x"0102", x"E030", x"24F8", x"7880", x"B9A0", x"7881",
   x"B9A1", x"0100", x"B9A2", x"B9A3", x"B9C0", x"B9C1", x"B9C2", x"B9C3",
   x"0101", x"E030", x"2505", x"7880", x"B9A0", x"0100", x"B9A1", x"B9A2",
   x"B9A3", x"B9C0", x"B9C1", x"B9C2", x"B9C3", x"7057", x"A053", x"B057",
   x"7802", x"2510", x"7058", x"A053", x"B058", x"7059", x"A053", x"B059",
   x"013B", x"B800", x"1526", x"678B", x"01EB", x"67C0", x"0128", x"67C0",
   x"67C3", x"0107", x"B800", x"66A0", x"1526", x"6759", x"0100", x"6705",
   x"3523", x"0108", x"B800", x"1526", x"1526", x"1526", x"7801", x"B980",
   x"7802", x"B981", x"7800", x"B982", x"780C", x"B983", x"0C20", x"0C90",
   x"0D01", x"0D84", x"7052", x"C052", x"B052", x"902A", x"B053", x"7044",
   x"E029", x"B044", x"205E", x"0110", x"E04C", x"254A", x"7055", x"902A",
   x"A04B", x"A057", x"B80C", x"A059", x"254A", x"7058", x"B402", x"0100",
   x"B04C", x"B400", x"0109", x"E04C", x"2556", x"7055", x"A056", x"A04B",
   x"2556", x"7055", x"B402", x"0100", x"B04C", x"B400", x"010F", x"E04C",
   x"2562", x"7055", x"A056", x"A04B", x"2562", x"7055", x"B402", x"0100",
   x"B04C", x"B400", x"1640", x"0100", x"B04D", x"7430", x"B03B", x"7431",
   x"B03C", x"7432", x"B03D", x"7433", x"B03E", x"01A0", x"B035", x"0186",
   x"B036", x"0101", x"B037", x"0100", x"B038", x"0100", x"B033", x"B034",
   x"0100", x"B039", x"B03A", x"66BC", x"7033", x"B422", x"7034", x"B423",
   x"0100", x"0980", x"0106", x"0B80", x"704A", x"C028", x"0200", x"0200",
   x"0200", x"B030", x"704A", x"C028", x"0200", x"0200", x"C030", x"B030",
   x"0001", x"0001", x"7030", x"B045", x"0100", x"B980", x"0D81", x"7045",
   x"E029", x"B045", x"2594", x"0180", x"0800", x"0100", x"0A00", x"0180",
   x"0900", x"0104", x"0B00", x"0100", x"0980", x"0106", x"0B80", x"0100",
   x"B04B", x"704A", x"B045", x"0100", x"B80B", x"B800", x"B801", x"B80C",
   x"01C1", x"B802", x"66A5", x"01A0", x"B033", x"0186", x"B034", x"0101",
   x"B035", x"0100", x"B036", x"0100", x"B037", x"0100", x"B038", x"0100",
   x"B039", x"0100", x"B03A", x"0164", x"B812", x"0100", x"B813", x"7818",
   x"B040", x"7819", x"B041", x"781A", x"B042", x"781B", x"B043", x"66AF",
   x"66AF", x"66AF", x"66AF", x"0100", x"B033", x"B034", x"B039", x"B03A",
   x"7040", x"B035", x"7041", x"B036", x"7042", x"B037", x"7043", x"B038",
   x"7430", x"B03B", x"7431", x"B03C", x"7432", x"B03D", x"7433", x"B03E",
   x"66BC", x"7034", x"260D", x"7037", x"C037", x"B037", x"7038", x"D038",
   x"B038", x"7039", x"D039", x"B039", x"703A", x"D03A", x"B03A", x"7037",
   x"E430", x"7038", x"F431", x"7039", x"F432", x"703A", x"F433", x"560C",
   x"0101", x"C033", x"B033", x"0100", x"D034", x"B034", x"0100", x"D035",
   x"B035", x"0100", x"D036", x"B036", x"1619", x"0101", x"C033", x"B033",
   x"0100", x"D034", x"B034", x"0100", x"D035", x"B035", x"0100", x"D036",
   x"B036", x"7033", x"B910", x"7034", x"B920", x"7035", x"B930", x"B940",
   x"0100", x"B950", x"0120", x"B970", x"7801", x"B980", x"7802", x"B981",
   x"7800", x"B982", x"780C", x"B983", x"01FF", x"C02A", x"704B", x"0200",
   x"B04B", x"0C20", x"0D01", x"0D84", x"7045", x"E029", x"B045", x"25AB",
   x"01FF", x"B049", x"0108", x"E401", x"2640", x"0100", x"B04C", x"B400",
   x"704C", x"264B", x"7401", x"364B", x"B02D", x"0A80", x"B04C", x"B04E",
   x"7400", x"B02C", x"0880", x"704E", x"369F", x"0120", x"A02D", x"365D",
   x"0100", x"B04E", x"0180", x"A02D", x"3658", x"7402", x"B880", x"165A",
   x"7880", x"B402", x"0100", x"B04C", x"B400", x"0110", x"A02D", x"3669",
   x"0100", x"B04E", x"702C", x"B057", x"B058", x"B059", x"01DE", x"A802",
   x"B802", x"704D", x"268D", x"0109", x"E02D", x"2680", x"01BD", x"B05C",
   x"7600", x"0101", x"E603", x"2676", x"01BF", x"B05C", x"0100", x"B04E",
   x"01FF", x"B04D", x"702D", x"B048", x"702C", x"B054", x"B055", x"B056",
   x"010F", x"E02D", x"268D", x"0100", x"B04E", x"01FF", x"B04D", x"702D",
   x"B048", x"702C", x"B054", x"B055", x"B056", x"0108", x"E02D", x"2698",
   x"0100", x"B04E", x"0100", x"B049", x"B04D", x"B054", x"B048", x"B402",
   x"704E", x"369F", x"0100", x"B04E", x"0100", x"B04C", x"B400", x"1046",
   x"7422", x"B810", x"7423", x"B811", x"1800", x"0100", x"B803", x"B804",
   x"B805", x"B806", x"B807", x"B808", x"01C8", x"B809", x"1800", x"7040",
   x"C040", x"B040", x"7041", x"D041", x"B041", x"7042", x"D042", x"B042",
   x"7043", x"D043", x"B043", x"1800", x"011F", x"B03F", x"7033", x"C033",
   x"B033", x"7034", x"D034", x"B034", x"7035", x"D035", x"B035", x"7036",
   x"D036", x"B036", x"7037", x"D037", x"B037", x"7038", x"D038", x"B038",
   x"7039", x"D039", x"B039", x"703A", x"D03A", x"B03A", x"56F5", x"7037",
   x"E03B", x"B037", x"7038", x"F03C", x"B038", x"7039", x"F03D", x"B039",
   x"703A", x"F03E", x"B03A", x"46F1", x"7037", x"C03B", x"B037", x"7038",
   x"D03C", x"B038", x"7039", x"D03D", x"B039", x"703A", x"D03E", x"B03A",
   x"16F4", x"0101", x"C033", x"B033", x"16FE", x"7037", x"E03B", x"B037",
   x"7038", x"F03C", x"B038", x"0101", x"C033", x"B033", x"703F", x"E029",
   x"B03F", x"46BE", x"0003", x"0003", x"1800", x"B02E", x"C029", x"B02F",
   x"B425", x"7940", x"E02F", x"5757", x"702E", x"3721", x"0480", x"B05A",
   x"0680", x"B05B", x"0003", x"0003", x"7900", x"B880", x"B424", x"0C81",
   x"702E", x"E029", x"B02E", x"2712", x"705A", x"0880", x"705B", x"0A80",
   x"0003", x"7900", x"E424", x"3754", x"0101", x"C803", x"572A", x"B803",
   x"0003", x"173F", x"7809", x"E803", x"473F", x"0180", x"8801", x"B801",
   x"7059", x"A053", x"B059", x"0180", x"A801", x"3739", x"7056", x"A053",
   x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"0101",
   x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"374B",
   x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100",
   x"B950", x"0180", x"0200", x"1755", x"C028", x"01FF", x"1758", x"0100",
   x"1800", x"7422", x"E810", x"E812", x"578A", x"0101", x"C806", x"5763",
   x"B806", x"0003", x"1778", x"7809", x"E806", x"4778", x"0180", x"8801",
   x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"3772", x"7056",
   x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950",
   x"0108", x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801",
   x"3784", x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940",
   x"0100", x"B950", x"1800", x"0003", x"7960", x"278B", x"B425", x"7940",
   x"37BF", x"0101", x"C807", x"5797", x"B807", x"0003", x"17AC", x"7809",
   x"E807", x"47AC", x"0180", x"8801", x"B801", x"7059", x"A053", x"B059",
   x"0180", x"A801", x"37A6", x"7056", x"A053", x"B056", x"0120", x"8802",
   x"B802", x"B940", x"0100", x"B950", x"0110", x"8801", x"B801", x"7059",
   x"A053", x"B059", x"0180", x"A801", x"37B8", x"7056", x"A053", x"B056",
   x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"B940", x"1800",
   x"B424", x"B900", x"1800", x"7424", x"B900", x"1800", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"ABCD"
);

signal daddra: std_logic_vector(10 downto 0);
signal daddrb: std_logic_vector(10 downto 0);

begin
   asslbp: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (wea = '1') then
            RAM(conv_integer(addra)) <= dina;
         end if;
         daddra <= addra;
         daddrb <= addrb;
      end if; -- clk 
   end process;

   douta <= RAM(conv_integer(daddra));
   doutb <= RAM(conv_integer(daddrb));
end;
