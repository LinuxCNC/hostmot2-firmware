library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from zero.bin
-- On12/31/2008

entity testram is
	port (
	addra: in std_logic_vector(10 downto 0);
	addrb: in std_logic_vector(10 downto 0);
	clk: in std_logic;
	dina: in std_logic_vector(31 downto 0);
	douta: out std_logic_vector(31 downto 0);
	doutb: out std_logic_vector(31 downto 0);
	wea: in std_logic);
end testram;

architecture syn of testram is
   type ram_type is array (0 to 2047) of std_logic_vector(31 downto 0);
   signal RAM : ram_type := 
   (
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000",
   x"00000000", x"00000000", x"00000000", x"00000000"
);

signal daddra: std_logic_vector(10 downto 0);
signal daddrb: std_logic_vector(10 downto 0);

begin
   atestram: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (wea = '1') then
            RAM(conv_integer(addra)) <= dina;
         end if;
         daddra <= addra;
         daddrb <= addrb;
      end if; -- clk 
   end process;

   douta <= RAM(conv_integer(daddra));
   doutb <= RAM(conv_integer(daddrb));
end;
