library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from sslbp.bin
-- On 12/15/2010

entity sslbp is
	port (
	addra: in std_logic_vector(10 downto 0);
	addrb: in std_logic_vector(10 downto 0);
	clk: in std_logic;
	dina: in std_logic_vector(15 downto 0);
	douta: out std_logic_vector(15 downto 0);
	doutb: out std_logic_vector(15 downto 0);
	wea: in std_logic);
end sslbp;

architecture syn of sslbp is
   type ram_type is array (0 to 2047) of std_logic_vector(15 downto 0);
   signal RAM : ram_type := 
   (
   x"0000", x"0000", x"0100", x"B028", x"B054", x"B049", x"B04C", x"0101",
   x"B029", x"01FF", x"B02A", x"0155", x"B02B", x"01AA", x"B402", x"7434",
   x"B04A", x"0138", x"B008", x"0149", x"B009", x"0132", x"B00A", x"0130",
   x"B00B", x"0137", x"B00C", x"0149", x"B00D", x"0136", x"B00E", x"0134",
   x"B00F", x"0112", x"B000", x"0101", x"B002", x"010D", x"B003", x"0108",
   x"B001", x"01D8", x"B006", x"704A", x"B007", x"0180", x"0800", x"0100",
   x"0A00", x"0002", x"704A", x"B045", x"01A0", x"B818", x"0125", x"B819",
   x"0126", x"B81A", x"0100", x"B81B", x"0C20", x"7045", x"E029", x"B045",
   x"2034", x"0100", x"B049", x"0100", x"B04C", x"B400", x"7049", x"355B",
   x"0180", x"0800", x"0100", x"0A00", x"0180", x"0880", x"0101", x"0A80",
   x"0180", x"0900", x"0104", x"0B00", x"0100", x"0980", x"0106", x"0B80",
   x"0101", x"B052", x"01FE", x"B053", x"704A", x"B044", x"0180", x"A801",
   x"251E", x"7054", x"A052", x"351E", x"016B", x"C800", x"0E80", x"0000",
   x"0000", x"0000", x"1800", x"11B3", x"11B8", x"11BC", x"11CA", x"11D2",
   x"11DD", x"150B", x"1515", x"1212", x"121C", x"1223", x"122B", x"1232",
   x"1237", x"123F", x"1246", x"1251", x"1259", x"1260", x"126A", x"1271",
   x"127B", x"1282", x"128C", x"1293", x"12BF", x"1305", x"1315", x"131C",
   x"1328", x"132F", x"1338", x"1344", x"134B", x"1386", x"1396", x"139D",
   x"13AD", x"13B4", x"13C0", x"13C7", x"13D0", x"13DC", x"13E3", x"1421",
   x"1431", x"10F1", x"10F9", x"1100", x"10AB", x"10C0", x"10CE", x"12EB",
   x"12FB", x"1189", x"1199", x"1142", x"1157", x"1165", x"143C", x"14B0",
   x"14BB", x"151C", x"151D", x"7057", x"A052", x"30BF", x"0003", x"0003",
   x"6772", x"705C", x"67A6", x"79A0", x"67A6", x"79A1", x"67A6", x"79A2",
   x"67A6", x"79A3", x"67A6", x"67A9", x"6689", x"0132", x"B800", x"151E",
   x"6741", x"50C4", x"0131", x"B800", x"0108", x"66EE", x"30CD", x"40CB",
   x"0131", x"B800", x"10CD", x"0133", x"B800", x"151E", x"7880", x"B9C0",
   x"7881", x"B9C1", x"7882", x"B9C2", x"7883", x"B9C3", x"8882", x"30DB",
   x"0101", x"8802", x"B802", x"7886", x"B9A0", x"7887", x"B9A1", x"7884",
   x"B9A2", x"7885", x"B9A3", x"7057", x"A053", x"B057", x"7802", x"20EE",
   x"7058", x"A053", x"B058", x"7059", x"A053", x"B059", x"0131", x"B800",
   x"151E", x"6772", x"01DF", x"67A6", x"67A9", x"012F", x"B800", x"6689",
   x"151E", x"6741", x"0101", x"66EE", x"30FF", x"0130", x"B800", x"151E",
   x"015A", x"E880", x"2115", x"017F", x"A802", x"B802", x"7055", x"A053",
   x"B055", x"7056", x"A053", x"B056", x"7057", x"A052", x"3112", x"0131",
   x"B800", x"1114", x"012E", x"B800", x"1141", x"7804", x"E809", x"411D",
   x"0101", x"C804", x"B804", x"0003", x"112F", x"0180", x"8801", x"B801",
   x"7059", x"A053", x"B059", x"0180", x"A801", x"3129", x"7056", x"A053",
   x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"0102",
   x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"313B",
   x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100",
   x"B950", x"151E", x"7057", x"A052", x"3156", x"0003", x"0003", x"6772",
   x"705C", x"67A6", x"79A0", x"67A6", x"79A1", x"67A6", x"79A2", x"67A6",
   x"0100", x"67A6", x"67A9", x"6689", x"0139", x"B800", x"151E", x"6741",
   x"515B", x"0138", x"B800", x"0108", x"66EE", x"3164", x"4162", x"0138",
   x"B800", x"1164", x"013A", x"B800", x"151E", x"7880", x"B9A0", x"7881",
   x"B9A1", x"7882", x"B9A2", x"0108", x"A883", x"3171", x"0101", x"8802",
   x"B802", x"0100", x"B9A3", x"7884", x"B9C0", x"7885", x"B9C1", x"7886",
   x"B9C2", x"7887", x"B9C3", x"7057", x"A053", x"B057", x"7802", x"2186",
   x"7058", x"A053", x"B058", x"7059", x"A053", x"B059", x"0138", x"B800",
   x"151E", x"6772", x"705C", x"67A6", x"0100", x"67A6", x"0100", x"67A6",
   x"0100", x"67A6", x"0100", x"67A6", x"67A9", x"0137", x"B800", x"6689",
   x"151E", x"6741", x"0108", x"66EE", x"31B2", x"017F", x"A802", x"B802",
   x"7055", x"A053", x"B055", x"7056", x"A053", x"B056", x"7057", x"A052",
   x"31AC", x"0138", x"B800", x"11B2", x"0128", x"B812", x"0100", x"B813",
   x"0136", x"B800", x"151E", x"668E", x"B940", x"0101", x"B800", x"151E",
   x"6689", x"0102", x"B800", x"151E", x"7422", x"E810", x"B031", x"7423",
   x"F811", x"B032", x"7812", x"E031", x"7813", x"F032", x"41C9", x"0103",
   x"B800", x"151E", x"6772", x"01DF", x"67A6", x"67A9", x"0104", x"B800",
   x"6689", x"151E", x"6741", x"51D7", x"0101", x"B800", x"11DC", x"0101",
   x"66EE", x"31DC", x"0105", x"B800", x"151E", x"015A", x"E880", x"21E3",
   x"0106", x"B800", x"1211", x"7804", x"E809", x"41EB", x"0101", x"C804",
   x"B804", x"0003", x"11FD", x"0180", x"8801", x"B801", x"7059", x"A053",
   x"B059", x"0180", x"A801", x"31F7", x"7056", x"A053", x"B056", x"0120",
   x"8802", x"B802", x"B940", x"0100", x"B950", x"0102", x"8801", x"B801",
   x"7059", x"A053", x"B059", x"0180", x"A801", x"3209", x"7056", x"A053",
   x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"0101",
   x"B800", x"151E", x"6772", x"01E1", x"67A6", x"0100", x"67A6", x"67A9",
   x"0109", x"B800", x"6689", x"151E", x"6741", x"0100", x"66EE", x"3222",
   x"010A", x"B800", x"151E", x"6772", x"01C1", x"67A6", x"67A9", x"010B",
   x"B800", x"6689", x"151E", x"6741", x"0101", x"66EE", x"3231", x"010C",
   x"B800", x"151E", x"7880", x"2236", x"010D", x"B800", x"151E", x"6772",
   x"01BC", x"67A6", x"67A9", x"010E", x"B800", x"6689", x"151E", x"6741",
   x"0104", x"66EE", x"3245", x"010F", x"B800", x"151E", x"7880", x"B9A0",
   x"7881", x"B9A1", x"7882", x"B9A2", x"7883", x"B9A3", x"0110", x"B800",
   x"151E", x"6772", x"01D0", x"67A6", x"67A9", x"0111", x"B800", x"6689",
   x"151E", x"6741", x"0101", x"66EE", x"325F", x"0112", x"B800", x"151E",
   x"7880", x"B814", x"6772", x"01D1", x"67A6", x"67A9", x"0113", x"B800",
   x"6689", x"151E", x"6741", x"0101", x"66EE", x"3270", x"0114", x"B800",
   x"151E", x"7880", x"B815", x"6772", x"01D2", x"67A6", x"67A9", x"0115",
   x"B800", x"6689", x"151E", x"6741", x"0101", x"66EE", x"3281", x"0116",
   x"B800", x"151E", x"7880", x"B816", x"6772", x"01D3", x"67A6", x"67A9",
   x"0117", x"B800", x"6689", x"151E", x"6741", x"0101", x"66EE", x"3292",
   x"0118", x"B800", x"151E", x"0119", x"B800", x"7880", x"B817", x"7008",
   x"E814", x"B030", x"7009", x"F815", x"8030", x"B030", x"700A", x"F816",
   x"8030", x"B030", x"700B", x"F817", x"8030", x"22BE", x"0180", x"B80C",
   x"0109", x"E048", x"22B0", x"01BF", x"A802", x"B802", x"011A", x"B800",
   x"010F", x"E048", x"22BE", x"013E", x"A802", x"B802", x"7055", x"A053",
   x"B055", x"7056", x"A053", x"B056", x"013B", x"B800", x"151E", x"013F",
   x"B800", x"7880", x"B817", x"700C", x"E814", x"B030", x"700D", x"F815",
   x"8030", x"B030", x"700E", x"F816", x"8030", x"B030", x"700F", x"F817",
   x"8030", x"22EA", x"0174", x"B80C", x"0109", x"E048", x"22DC", x"01BF",
   x"A802", x"B802", x"0134", x"B800", x"010F", x"E048", x"22EA", x"013E",
   x"A802", x"B802", x"7055", x"A053", x"B055", x"7056", x"A053", x"B056",
   x"013B", x"B800", x"151E", x"6772", x"705C", x"67A6", x"0100", x"67A6",
   x"0100", x"67A6", x"0100", x"67A6", x"0108", x"67A6", x"67A9", x"0135",
   x"B800", x"6689", x"151E", x"6741", x"0108", x"66EE", x"3304", x"01FE",
   x"A802", x"B802", x"0136", x"B800", x"151E", x"6772", x"0165", x"67A6",
   x"0154", x"67A6", x"0108", x"67A6", x"01FF", x"67A6", x"01FF", x"67A6",
   x"67A9", x"011B", x"B800", x"6689", x"151E", x"6741", x"0100", x"66EE",
   x"331B", x"011C", x"B800", x"151E", x"6772", x"0145", x"67A6", x"0154",
   x"67A6", x"0108", x"67A6", x"67A9", x"011D", x"B800", x"6689", x"151E",
   x"6741", x"0102", x"66EE", x"332E", x"011E", x"B800", x"151E", x"7880",
   x"8881", x"2335", x"011F", x"B800", x"1337", x"011C", x"B800", x"151E",
   x"6772", x"0145", x"67A6", x"0152", x"67A6", x"0108", x"67A6", x"67A9",
   x"0120", x"B800", x"6689", x"151E", x"6741", x"0102", x"66EE", x"334A",
   x"0121", x"B800", x"151E", x"0180", x"B9C0", x"0100", x"B9C1", x"7880",
   x"B9C2", x"7881", x"B9C3", x"7880", x"8881", x"2359", x"0122", x"B800",
   x"1385", x"7808", x"E809", x"4361", x"0101", x"C808", x"B808", x"0003",
   x"1373", x"0180", x"8801", x"B801", x"7059", x"A053", x"B059", x"0180",
   x"A801", x"336D", x"7056", x"A053", x"B056", x"0120", x"8802", x"B802",
   x"B940", x"0100", x"B950", x"0140", x"8801", x"B801", x"7059", x"A053",
   x"B059", x"0180", x"A801", x"337F", x"7056", x"A053", x"B056", x"0120",
   x"8802", x"B802", x"B940", x"0100", x"B950", x"151E", x"6772", x"0165",
   x"67A6", x"0160", x"67A6", x"0108", x"67A6", x"0100", x"67A6", x"0100",
   x"67A6", x"67A9", x"0123", x"B800", x"6689", x"151E", x"6741", x"0100",
   x"66EE", x"339C", x"0124", x"B800", x"151E", x"6772", x"0165", x"67A6",
   x"0104", x"67A6", x"0108", x"67A6", x"01FF", x"67A6", x"01FF", x"67A6",
   x"67A9", x"0125", x"B800", x"6689", x"151E", x"6741", x"0100", x"66EE",
   x"33B3", x"0126", x"B800", x"151E", x"6772", x"0145", x"67A6", x"01FE",
   x"67A6", x"0108", x"67A6", x"67A9", x"0127", x"B800", x"6689", x"151E",
   x"6741", x"0102", x"66EE", x"33C6", x"0128", x"B800", x"151E", x"7880",
   x"8881", x"23CD", x"0126", x"B800", x"13CF", x"0129", x"B800", x"151E",
   x"6772", x"0145", x"67A6", x"0152", x"67A6", x"0108", x"67A6", x"67A9",
   x"012A", x"B800", x"6689", x"151E", x"6741", x"0102", x"66EE", x"33E2",
   x"012B", x"B800", x"151E", x"0180", x"B9C0", x"0100", x"B9C1", x"7880",
   x"B9C2", x"7881", x"B9C3", x"7880", x"8881", x"23F4", x"01FE", x"A802",
   x"B802", x"012C", x"B800", x"1420", x"7808", x"E809", x"43FC", x"0101",
   x"C808", x"B808", x"0003", x"140E", x"0180", x"8801", x"B801", x"7059",
   x"A053", x"B059", x"0180", x"A801", x"3408", x"7056", x"A053", x"B056",
   x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"0140", x"8801",
   x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"341A", x"7056",
   x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950",
   x"151E", x"6772", x"0165", x"67A6", x"015C", x"67A6", x"0108", x"67A6",
   x"01F4", x"67A6", x"0101", x"67A6", x"67A9", x"012D", x"B800", x"6689",
   x"151E", x"6741", x"0100", x"66EE", x"343B", x"010F", x"B812", x"0100",
   x"B813", x"012E", x"B800", x"151E", x"0164", x"B812", x"0100", x"B813",
   x"7057", x"A052", x"34AF", x"0003", x"0003", x"6772", x"7980", x"B050",
   x"7981", x"B051", x"7983", x"B04F", x"67A6", x"0103", x"A04F", x"B046",
   x"C028", x"0101", x"B047", x"7046", x"345E", x"7047", x"0200", x"B047",
   x"7046", x"E029", x"B046", x"0001", x"0001", x"1453", x"01BF", x"E04F",
   x"54A0", x"0104", x"A04F", x"3469", x"0003", x"7050", x"67A6", x"7051",
   x"67A6", x"0120", x"A04F", x"349D", x"0100", x"B80A", x"0108", x"E047",
   x"2482", x"0003", x"79A0", x"67A6", x"79A1", x"67A6", x"79A2", x"67A6",
   x"79A3", x"67A6", x"79C0", x"67A6", x"79C1", x"67A6", x"79C2", x"67A6",
   x"79C3", x"67A6", x"0104", x"E047", x"248E", x"0003", x"79A0", x"67A6",
   x"79A1", x"67A6", x"79A2", x"67A6", x"79A3", x"67A6", x"0102", x"E047",
   x"2496", x"0003", x"79A0", x"67A6", x"79A1", x"67A6", x"0101", x"E047",
   x"249C", x"0003", x"79A0", x"67A6", x"149F", x"7047", x"B80A", x"14AB",
   x"0120", x"A04F", x"34A9", x"0003", x"79A0", x"67A6", x"0100", x"B80A",
   x"14AB", x"0101", x"B80A", x"67A9", x"6689", x"013C", x"B800", x"151E",
   x"6741", x"780A", x"66EE", x"34BA", x"44B8", x"013B", x"B800", x"14BA",
   x"013D", x"B800", x"151E", x"780A", x"B030", x"0001", x"0001", x"0108",
   x"E030", x"24D2", x"7880", x"B9A0", x"7881", x"B9A1", x"7882", x"B9A2",
   x"7883", x"B9A3", x"7884", x"B9C0", x"7885", x"B9C1", x"7886", x"B9C2",
   x"7887", x"B9C3", x"0104", x"E030", x"24E2", x"7880", x"B9A0", x"7881",
   x"B9A1", x"7882", x"B9A2", x"7883", x"B9A3", x"0100", x"B9C0", x"B9C1",
   x"B9C2", x"B9C3", x"0102", x"E030", x"24F0", x"7880", x"B9A0", x"7881",
   x"B9A1", x"0100", x"B9A2", x"B9A3", x"B9C0", x"B9C1", x"B9C2", x"B9C3",
   x"0101", x"E030", x"24FD", x"7880", x"B9A0", x"0100", x"B9A1", x"B9A2",
   x"B9A3", x"B9C0", x"B9C1", x"B9C2", x"B9C3", x"7057", x"A053", x"B057",
   x"7802", x"2508", x"7058", x"A053", x"B058", x"7059", x"A053", x"B059",
   x"013B", x"B800", x"151E", x"6772", x"01EB", x"67A6", x"0128", x"67A6",
   x"67A9", x"0107", x"B800", x"6689", x"151E", x"6741", x"0100", x"66EE",
   x"351B", x"0108", x"B800", x"151E", x"151E", x"151E", x"7801", x"B980",
   x"7802", x"B981", x"7800", x"B982", x"780C", x"B983", x"0C20", x"0C90",
   x"0D01", x"0D84", x"7052", x"C052", x"B052", x"902A", x"B053", x"7044",
   x"E029", x"B044", x"205E", x"0110", x"E04C", x"2542", x"7055", x"902A",
   x"A04B", x"A057", x"B80C", x"A059", x"2542", x"7058", x"B402", x"0100",
   x"B04C", x"B400", x"0109", x"E04C", x"254E", x"7055", x"A056", x"A04B",
   x"254E", x"7055", x"B402", x"0100", x"B04C", x"B400", x"010F", x"E04C",
   x"255A", x"7055", x"A056", x"A04B", x"255A", x"7055", x"B402", x"0100",
   x"B04C", x"B400", x"1611", x"0100", x"B04D", x"0100", x"0980", x"0106",
   x"0B80", x"015F", x"B045", x"0100", x"B980", x"0D81", x"7045", x"E029",
   x"B045", x"4563", x"0180", x"0800", x"0100", x"0A00", x"0180", x"0900",
   x"0104", x"0B00", x"0100", x"0980", x"0106", x"0B80", x"0100", x"B04B",
   x"704A", x"B045", x"0100", x"B80B", x"B800", x"B801", x"B80C", x"0114",
   x"B809", x"01C1", x"B802", x"668E", x"01A0", x"B033", x"0186", x"B034",
   x"0101", x"B035", x"0100", x"B036", x"0100", x"B037", x"0100", x"B038",
   x"0100", x"B039", x"0100", x"B03A", x"0164", x"B812", x"0100", x"B813",
   x"7818", x"B040", x"7819", x"B041", x"781A", x"B042", x"781B", x"B043",
   x"6698", x"6698", x"6698", x"6698", x"0100", x"B033", x"B034", x"B039",
   x"B03A", x"7040", x"B035", x"7041", x"B036", x"7042", x"B037", x"7043",
   x"B038", x"7430", x"B03B", x"7431", x"B03C", x"7432", x"B03D", x"7433",
   x"B03E", x"66A5", x"7034", x"25DE", x"7037", x"C037", x"B037", x"7038",
   x"D038", x"B038", x"7039", x"D039", x"B039", x"703A", x"D03A", x"B03A",
   x"7037", x"E430", x"7038", x"F431", x"7039", x"F432", x"703A", x"F433",
   x"55DD", x"0101", x"C033", x"B033", x"0100", x"D034", x"B034", x"0100",
   x"D035", x"B035", x"0100", x"D036", x"B036", x"15EA", x"0101", x"C033",
   x"B033", x"0100", x"D034", x"B034", x"0100", x"D035", x"B035", x"0100",
   x"D036", x"B036", x"7033", x"B910", x"7034", x"B920", x"7035", x"B930",
   x"B940", x"0100", x"B950", x"0120", x"B970", x"7801", x"B980", x"7802",
   x"B981", x"7800", x"B982", x"780C", x"B983", x"01FF", x"C02A", x"704B",
   x"0200", x"B04B", x"0C20", x"0D01", x"0D84", x"7045", x"E029", x"B045",
   x"257A", x"01FF", x"B049", x"0108", x"E401", x"2611", x"0100", x"B04C",
   x"B400", x"704C", x"261C", x"7401", x"361C", x"B02D", x"0A80", x"B04C",
   x"B04E", x"7400", x"B02C", x"0880", x"704E", x"3688", x"0120", x"A02D",
   x"362E", x"0100", x"B04E", x"0180", x"A02D", x"3629", x"7402", x"B880",
   x"162B", x"7880", x"B402", x"0100", x"B04C", x"B400", x"0110", x"A02D",
   x"3640", x"704D", x"363D", x"0100", x"B04E", x"702C", x"B057", x"B058",
   x"B059", x"01DE", x"A802", x"B802", x"1640", x"0100", x"B04C", x"B400",
   x"704D", x"2676", x"0109", x"E02D", x"2660", x"01A0", x"B05D", x"0186",
   x"B05E", x"0101", x"B05F", x"0100", x"B060", x"67AC", x"01BD", x"B05C",
   x"7600", x"0101", x"E603", x"2656", x"01BF", x"B05C", x"0100", x"B04E",
   x"01FF", x"B04D", x"702D", x"B048", x"702C", x"B054", x"B055", x"B056",
   x"010F", x"E02D", x"2676", x"01D0", x"B05D", x"0107", x"B05E", x"0100",
   x"B05F", x"0100", x"B060", x"67AC", x"0100", x"B04E", x"01FF", x"B04D",
   x"702D", x"B048", x"702C", x"B054", x"B055", x"B056", x"0108", x"E02D",
   x"2681", x"0100", x"B04E", x"0100", x"B049", x"B04D", x"B054", x"B048",
   x"B402", x"704E", x"3688", x"0100", x"B04E", x"0100", x"B04C", x"B400",
   x"1046", x"7422", x"B810", x"7423", x"B811", x"1800", x"0100", x"B803",
   x"B804", x"B805", x"B806", x"B807", x"B808", x"0114", x"B809", x"1800",
   x"7040", x"C040", x"B040", x"7041", x"D041", x"B041", x"7042", x"D042",
   x"B042", x"7043", x"D043", x"B043", x"1800", x"011F", x"B03F", x"7033",
   x"C033", x"B033", x"7034", x"D034", x"B034", x"7035", x"D035", x"B035",
   x"7036", x"D036", x"B036", x"7037", x"D037", x"B037", x"7038", x"D038",
   x"B038", x"7039", x"D039", x"B039", x"703A", x"D03A", x"B03A", x"56DE",
   x"7037", x"E03B", x"B037", x"7038", x"F03C", x"B038", x"7039", x"F03D",
   x"B039", x"703A", x"F03E", x"B03A", x"46DA", x"7037", x"C03B", x"B037",
   x"7038", x"D03C", x"B038", x"7039", x"D03D", x"B039", x"703A", x"D03E",
   x"B03A", x"16DD", x"0101", x"C033", x"B033", x"16E7", x"7037", x"E03B",
   x"B037", x"7038", x"F03C", x"B038", x"0101", x"C033", x"B033", x"703F",
   x"E029", x"B03F", x"46A7", x"0003", x"0003", x"1800", x"B02E", x"C029",
   x"B02F", x"B425", x"7940", x"E02F", x"573F", x"702E", x"370A", x"0480",
   x"B05A", x"0680", x"B05B", x"0003", x"0003", x"7900", x"B880", x"B424",
   x"0C81", x"702E", x"E029", x"B02E", x"26FB", x"705A", x"0880", x"705B",
   x"0A80", x"0003", x"7900", x"E424", x"373C", x"7803", x"E809", x"4715",
   x"0101", x"C803", x"B803", x"0003", x"1727", x"0180", x"8801", x"B801",
   x"7059", x"A053", x"B059", x"0180", x"A801", x"3721", x"7056", x"A053",
   x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"0101",
   x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"3733",
   x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100",
   x"B950", x"0180", x"0200", x"173D", x"C028", x"01FF", x"1740", x"0100",
   x"1800", x"7422", x"E810", x"E812", x"5771", x"7806", x"E809", x"474D",
   x"0101", x"C806", x"B806", x"0003", x"175F", x"0180", x"8801", x"B801",
   x"7059", x"A053", x"B059", x"0180", x"A801", x"3759", x"7056", x"A053",
   x"B056", x"0120", x"8802", x"B802", x"B940", x"0100", x"B950", x"0108",
   x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801", x"376B",
   x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940", x"0100",
   x"B950", x"1800", x"0003", x"7960", x"2772", x"B425", x"7940", x"37A5",
   x"7807", x"E809", x"4780", x"0101", x"C807", x"B807", x"0003", x"1792",
   x"0180", x"8801", x"B801", x"7059", x"A053", x"B059", x"0180", x"A801",
   x"378C", x"7056", x"A053", x"B056", x"0120", x"8802", x"B802", x"B940",
   x"0100", x"B950", x"0110", x"8801", x"B801", x"7059", x"A053", x"B059",
   x"0180", x"A801", x"379E", x"7056", x"A053", x"B056", x"0120", x"8802",
   x"B802", x"B940", x"0100", x"B950", x"B940", x"1800", x"B424", x"B900",
   x"1800", x"7424", x"B900", x"1800", x"0E00", x"7430", x"B033", x"7431",
   x"B034", x"7432", x"B035", x"7433", x"B036", x"705D", x"B03B", x"705E",
   x"B03C", x"705F", x"B03D", x"7060", x"B03E", x"0100", x"B037", x"B038",
   x"0100", x"B039", x"B03A", x"66A5", x"0F00", x"7033", x"B061", x"7034",
   x"B062", x"7061", x"E029", x"B061", x"7062", x"F028", x"B062", x"7061",
   x"E029", x"B061", x"7062", x"F028", x"B062", x"7061", x"B422", x"7062",
   x"B423", x"1800", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"ABCD"
);

signal daddra: std_logic_vector(10 downto 0);
signal daddrb: std_logic_vector(10 downto 0);

begin
   asslbp: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (wea = '1') then
            RAM(conv_integer(addra)) <= dina;
         end if;
         daddra <= addra;
         daddrb <= addrb;
      end if; -- clk 
   end process;

   douta <= RAM(conv_integer(daddra));
   doutb <= RAM(conv_integer(daddrb));
end;
